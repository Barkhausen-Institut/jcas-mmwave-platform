-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��G<�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mώ�0����S��C�����u�u�0�!�:�8�W��L���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�6�w�m�Bϝ�	����[��V������&�'�8�9�.�4�������\ǶN��ʇ�2�!�u�0�2�+���Y����\��'�����0�!�u�;�2�3�ϗ�����G��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z�p�W���	����9K�c��U���%�;�;�u�9�)��������"��V����:�;�u�;�w�<�Ϫ�Ӕ��F
��U��U���x�u�=�u�;�*����ӂ��R��'�����0�<�;�1�#�}�Ͻ�����Q
��@��U���u�c�_�x�6�9�$�������9K��C�����:�&�4�!�w�����Ӈ����C��"���=�6�;�7�w�.�Ϫ�Y����Z ��@��ʡ�0�x�u�:�3�3�W������/��RN�����0�!�1�!�>�}����������U�����&�_�x�x�w�<����Y���R��Z�����0�y�a�u�>�.�W������V��^������u�u�u�w�r�[��H����Z��SB��Dʷ�!�y�d�u�9�8�������K����9���o�u�w�e�g�m�G���?��ƴF��B�����!�u�h�f�l�p�}��-����\��_����u�'�u�0�9�}�����ƣ�UF��C��Uȧ� �1�:�!�6�9�UϬ�����l�:��ʼ�u�6�:�%�>�5�ϼ�Y����Z��vT�����3�&�u�:�/�m�G��I�Ɗ�u ǶN��[���d�u��&�6�8�P���Y����@��^ �����6�'�,�<�w�2�	������O�CחXʜ�u�=�u�:�9�}��������]F�@�U���;�!�0�;�:�8�W���	����Z����U��� �!�<�_�z�/����ӓ����YN����� �7�'�<�w�8����Ӓ����B�����:�;�0�u�8�3�Wϊ������[N�����<�u�u�0�8�?�����ƿ�T��DN�����'�u�9�0�3�}��������WH�c�����"�9�y�=� �+��������F��VN�����8�9�u�4�9�8����Yӯ��J	��E�����'� �1�;�]�p����Ӏ����DB�����=� �1� �2�)��������[�������;��7�� �4�������$�������'�u�:�;�>�:��������Q��F�����u�|�!�0�w�5�W�������\��Qd�U���!�;�u�{�w��W�������T	����U���;�u�;�u�?�}����������E�����e�_�x��#�.��������\��^ �����d�u�<�&�w�3�W���Y������X�����0�'�,�e�w�	����T�ƻ�@F��X��Dʙ��:�u�4�9�8��������U��^�U���;�&�_�x�z�}�W��+����~N��C�!���u�&�"�4�w�)�Ͻ�����Z��X���߇x�x�u�u�j��5���:����r4��~ חXʖ�i�u��9��?�}��8ɤ�F��C���������k�}�3���0����nl�=C����;�;�&�1�6�9��������@��V�����<�!�;�0�w�2����
����]F��RN��%�߇x�3�;�!�8�q��������AF�������u�:�u�:�4�3�W���Y����A��C��ʻ�4�u�4�=�]�p����Ӏ����^ �����:�0�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l��U��ʼ�0�n�u� �2�4��������T��_�[���n�u� �0�>�8�Y�������@��V�����u�,�!�0�>�}��������\ ��[����� ���n�"�8�"���0�Ț�\��Y��Ĕ��_�x�&�9�5��������_��h����!�!�u�$��-�����ƥ�9F��R �����u�u�>�<�2�8����Y�ƥ�G��EN�����g�!�u�u�j�o�^�ԜY����l�N�����u�u�u�u�w�3��������l�N�����;�u�u�u�w�3��������l��C��A���:�;�:�e�l�}�WϽ�����GF�N����&�1�9�2�4�+����Q����\��XN�N���u�6�6�;�9�.����Y����G��X	��*���!�'�g�u�8�3���B�����x�����1�o�:�!�$�9��������G	��W�����:�e�u�n�2�9�2���
����]��dװ���<�0�!�'�w�	�W���<����C4��Y
��U���_�u�:�%�9�3�W���M˃ƹF��R �����u�u�u����2���Y���F�N�����'�o�u�n�w�}�Wϟ�,����a#��N��U���o�<�!�2�%�g�W��Y���'��pN��U���u�u�u�u�m�4�������]ǻN��U������
��	�%���<����F�N��Oʷ�:�0�;�o�w��$��Y���'��x<��0������
���#���-����	F��E��U��w���w�]�}�W���&����gF�N��U���u�u�!�<�0�g�W͚�+����l�N��7�����u�u�w�}�W���Y����T��S��N���u�u���w�}�W���Y���F��^ �����o�u�n�u�w�}�5���)���F�N��U��&�'�;�u�j��>���-��ƹF�-��'�����u�u�w�}�MϷ�����\�UךU���u������2���Y�����R	��U��d�_�u�u�w��0���Y���F�N��U���0�0�u�h�f�W�W���Y����F�N��U���u�u�u�<��8����C�Ɣ�  ��q(��3���w�_�u�u�w��0���Y���F�N��U���0�0�u�h�f�W�W���Y����p'��n'��0���u�u�u�;�2�8�W��H���F�x>��1����u�u�u�w�}�W�������	[�d��U�������w�}�W���Y����Q��A�����h��e�e�g�m�G��[���F�g<��U���u�u�u�u�w�}�W�������	[�d��U�������w�}�W���Y����@��Y	��H�����n�u�w�}�$���)����a(�N��U��&�'�;�u�j��6���+����F�N��9��� ���
���W�������\�=��*����n�u�u�w��:���=���F�N��Oʦ�'�;�u�h�u��2��Y���3��h#��!���u�u�u�u�m�.����Y���~3��h=�����u�u��
��	�%���<����\��C����u��
���	�L���Y����`#��~#��U���u�u�u�o�$�/����D�ă�vR��UךU���:�!�_�u�w�}�;���Y���F�T�����!�
�9�2�4�W�W���Y���F�N��U���u�;�u�!��2��������T��S�����|�_�u�u�w��9���Y���F���U���
�:�<�
�2�)���Y����G	�UךU���u�� �u�w�}�W���CӉ����h�����0�!�'�g�w�2����I��ƹF�,��U���u�u�u�u�m�4�Wϭ�����Z��R����u�:�;�:�g�f�W���YӤ��}F�N��U���o�<�u�&�3�1��������AN��
�����e�n�u�u�w��8���Y���F�N��ʦ�1�9�2�6�!�>����Nӂ��]��G�U���u��u�u�w�}�W���Y�ƥ�F��S1�����#�6�:�}�`�9� ���Y����F�N��U���u�u�u�u�w�}��������T��A�����b�1�"�!�w�t�}���Y�Ɯ�z(�N��U���u�u�;�u�#�����&����\� N�����u�|�_�u�w�}�4���Y���F�T�� ���!�
�:�<��8����M�ƨ�D��^����u�u����}�W���Y����]F��C
�����6�_�u�u�w��%���-���F���U���
�:�<�
�2�)�������\F��d��U���������W���Y���@��B����u�u�u����6���,���	F��CN�����:�<�n�u�w�}�8���=���F�N����&�1�9�2�4�+����Q�ƨ�D��^����u�u����}�W���Y����]F��C
�����
�0�!�'�d�9� ���Y����F�N��'�����u�u�w�}��������T��A�����u�:�;�:�g�f�W���Yӫ��g5��y'��U���o�<�u�!��1����s���F��{:��2����u�u�u�"�}��������l�N��:�����u�u�w�}�W���Y����F
��^�U���u� ����
�W���Y�ƣ�GF��S1�����n�u�u�u��	�2���=����gF��X����� �:�<�n�w�}�Wώ�-����w#��t:��Oʺ�!�&�1� �8�4�L���Y����v'��N��U���u�o�<�u�$�9������ƹF�-��G���u�u�u�u�m�4�Wϭ�����T��=N��U�������w�}�W������G��[���ߊu�u�u��f�}�W���Y�������*���2�6�_�u�w�}�2��Y���F�T�����!�
�9�2�4�W�W���Y����F�N��U���u�;�u�!��1����s���F��t/��,���u�u�u�u�9�}��������l�N��6����u�u�u�w�}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u���;���+����F��^ ����� �:�<�n�w�}�Wϝ�)���F�N��Oʼ�u�&�1� �8�4�L���Y����`2��N��U���u�o�<�u�$�9������ƹF�<��4������u�m�4�Wϭ�����T��=N��U����� ���}�W������G��[���ߊu�u�u���}�W���Y�������*���2�6�_�u�w�}�$���Y���F�T�����!�
�9�2�4�W�W���Y����g4��N��U���u�;�u�!��1����s���F��c#��U���u�u�u�u�9�}��������l�N��'���u�u�u�u�w�}�W���Y����F
��^����;�u�:�%�9�3�L�ԜY����R
��g�����u�u�u�o�$�9��������G	��Y�����:�e�u�h��)����G���l�D������'�,�;�w�}�W��
����\��T��R��_�u�<�;�;�>����0����F�N�����2�6�o�u�g�f�}�������]��y��7���&�u�o�<�#�:���Y����V"��V��U��u�6�;�!�9�}�?���5���F���*���<�
�0�!�%�i�W������F��6��E��e�e���l�}��������X)��G�����u�u�;�0�2�}�J��B���T��=N��Xʁ�0�6�'�,�>�}��������R��N��Yʦ�u�1�u�;�#�8�W����ƿ�Z��[��ʼ�_�u�x�!�2��5ϭ�����[��C��3���u�u��'�.�3���s�Ƽ�\��DF���ߊu�0�<�_�w�}�Ϭ�
����V��-��\ʡ�0�_�u�u�w���������[��X��1����}�b�n�w�}������ƹ�������n�_�u��%�$���Y����A��e�����u��8��2�.�Eϻ�
�Ƣ�GF��V����|�_�_�&�c�8�������Vl��Y��ʸ�%�_�u�u�4�.����D�Ƨ�F��E��Y���u�u�'�g��}����Y����_��S����u�y�u�u�6�8�W�������q��DB��U���x�d�:�u�w��%���s���R��E�����!�0�;�1�#�>�W�������l�N�����&�!�%�!�2�3��������G��S�W����w�_�u�w�����Y���w/��t:�����u�6�&�'�0�`�W�������T�C��U���g��u�0�$�}�Wϼ������Z/�����u�u�u�x�f�2�W���;Ӵ��@l�N�����!�h�u����U�ԜY�Ư�A��Y��U��d�u�u�u�w�p�W���8����z(��r)ךU���4�'�<�&�;�8�W���I���F��R	��K��u�u�u�u�w�}�W��Y�Ə�a#��N�����u�k�-�f���1���?����F�Z��U��e�_�u�u�"�)��������[�BךU���%�:�0�0�w�c�G�ԜY�Ƽ�G��YN��U���e�e�e�e�g�m�[���YӖ��TF�_�U���u�u�u�u�w�p�Fώ�+��ƹF��R�����<�2�8�&�w�c�U���&����JǻN�����4�>�h�u���U�ԜY�ƿ�_9��C����u�����q�W�������F
��
P��;���w�_�u�u�$���������G��S�W������w�]�}�W���&����[�!��A���_�:�!�8�'�W�W������%��d��Uʴ�h�u��!��u�@Ϻ�����^�=N��U���k�6�4�4�9�l�W������JǻN��U��>�4�3�&�{�}�WϽ�����[�T-�����y�u�u�4�>�}�IϽ�����F��d��Uʷ�<�u�k�}�#�8���Y���l�N�����k�}�!�0�$�`�W��P���F��E�����;�h�u�e�{�}�Wϳ�����]��
P��E���u�u�4�:�#�`�W���6����F��d��Uʷ�:�!�h�u�'�3�}���Y����J��T��U��:�0�y�u�w�0��������[�X��Y���u�%�h�u��(��ԜY�Ƽ�G��Y�����u�k�:�0�{�}�WϮ�����W��T��Kʺ�0�y�u�u�8�8����Y����C��=N��U���0�3�:�u�i�2���Y����R��X��H���%�;�_�u�w�>����GӉ��]JǻN�����0�h�u�e�f�m�F��Y����_��S��K���e�e�y�u�w�>��������X�^�Y���u�6�4�u�i�z�P�ԜY�Ư�RT�	N��R�ߊu�u�0�9�:�9�W���^����F�T��U��r�r�_�u�w�8�E��Y���9F���U��r�r�_�u�w�8�������A��d��Uʶ�8�h�u�d�{�}�WϽ�����X�I�U���6�%�h�u�f�q�W�������G��E��U��r�r�_�u�w�.���Y���9F������:�0�h�u�g�q�W�������X�I�U���'�!�u�k�p�z�}���Y����_
��E����u�e�y�u�w�/����G����l�N�����9�h�u�e�{�}�WϬ����A��UװU���u�=�u��$�5��������\��R
�����>�0�u�=�w���������|��S��%���9�a�u�:�9�2�C���6����G1��C���1���_