-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��C��&���9�;�{�=�]�p�6�������R��V������<�<�4�w�/����CӶ��V9��OחXʑ�!�o�d��'�8����K����KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��t�E��Y����A��CN�����4�u�;�!�"�8��������R��Yd�U���u�<�=�&��.����s����R��Y��<���'�8�;�&��)����Y����A��^��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��)����@��C�����6�8�:�0�#�4��������G��Q��ʴ�1�'�4�1�$�?�����ƪ�AF��RN�����_�x�3�9�2�}��������F����ʧ� �1�u�=�w�����0�Ƹ�X��^ �����<�u�=�_�z�����:������V�����%�&�0�u�#�)�W���Y����_��\N�����{�u�=�u�9�(�W������Z��E�����&�6�u�=�#�u�^Ϸ�Y����]��D�����u��0�:�#�(�W���ӏ��R��Y	�����&�6�u�=�#�u�^Ϸ�Y����\
��D�����u��<�u�6�>�����ƀ� ��vN�����0�!�!�:�]�p����(ӂ��RHǶd�U���u��a�r�w�.�ϸ�Ӓ����R�����&�7�'�6�8�.��������WF�������u�=�_�x���Oȭ�����U	��C�����1�;�y�4�3�<�����Ƹ�VF��X�����<�6�:�&�9�s�W���
���Z��E�����3�'�8�0�>�:�����ƪ�\��_�����u�-�!�4�$�)���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�<�'�'�w�8��ԜY����Z����*���<�
�d�a�6�1�}���
�ƥ�V��B�����!�{�9�n�w�(�ϩ��Ȝ�T#��V�����4�9�_�0�#�)�W���6����G5��G�����2�0�<�_�w�8����Q�����TN��U���u�u�u�o�>�)��������T��XN�U��m�|�_�u�8�)�}���Y����_��\N��U���u�u�;�&�3�1����s���`��[��ح�u�u�u�u�9�.��������F�T<�����!�u�u�u�w�}�ϭ�����Z��=N��U���!��u�u�w�}�W���Ɵ�P"��V1��]���6�g�x�u�8�3���B�����C�����;�u�u�o�>�}��������9l�N����� �u�u�u�w�}�W���Y����F��C��]���6�d�1�"�#�}�^�ԶY����w��a�����u�u�o�:�#�.�������l��SN�����%�!�4�%�>�:������ƓR��^�����u��u�3��-��������_��d�����&�_�u�x�?�2�(���
����9F������<�0�1�_�w�4��������z��NN��U����!�
�}�<�-�X���Hӂ��]��G��H���!�0�&�k�8�5���^���l�D������!���"�9����Cӵ��w��h��&���d�1�"�!�w�t�M�������@[�X����r�r�|�_�w�$����8����P��h��ʴ�'�,�}�;�2�8�W������	��D�����6�#�6�:��d��������l�D������!��9�3�2����Cӕ��l
��^�����'�f�1�"�#�}�^��Yۉ��V��	I�\�ߠ7�2�;�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F�/�����4�1��7�%�>��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�U���u�&�&���e�Ϫ�Y����F��T*������x�6�4�6�3�4���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�'�4�2�1��ԜY����V��d�����>�-�_�u�2�4�}���Y����Z��P1�����4�%�0�9�e�t����s���F��V�����u�h�6�4�6�3�}���Y����Z ��N��ʥ�:�0�&�_�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�����0�&�u�:�w�+�ϰ�����\ ��X�����;�&�u�x�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�������m�&�#�}����Y����zF��SN�����{�u�=�&�$�>��������^	��DN��ʱ�!�_�u�x�5�>�W�������R��R-��U���4�;�u��2�.��������GF����ʳ�'�0�0�u�w�9�}���Tӈ��Q��X�����<�<�;�&�2�-����Y����G�������0�1�3�0�2�>�W�������P��=N��Xʳ�'� �&�'�6�s�W��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠu�x�u�0�?�-�W�������A	��D��1�����,�u��)�>���T����R'��d��\���7�2�;�u�w�p�W��Y���O��^��Eʓ�&�u�u�6�6�<��������V�S��1����}�|�_�w�}�Z���P���U�@��U����u�u�x�w�o�W��Q����Z��N�����u�x�}�|�k�}�F������ ��N��X���a�u�h�}�~�*����Y��ƹF��X��U���d�!�u��4�o����s���F��V�����;�0���w�`��������JN��d��G���|�_�u�u�9�}����s���K�G��H���|�"�!�u�w��W���T���F�F�U���=�e��_�w�}�Z���P���W�@��U����u�u�3�%���������O������x�u�:�%�w�}�WϽ�����a	��S��]���i�u��!��u�$���0��ƹF��Y
�����_�u�;�u�%�>���s�Ƌ�]4��Y
���ߊu�:�u�u�9�m����*�����R���ߊu�u�0�f�>�8�}���Y����V��R �����_�u�u�u�z�5����Y����@��B ��ʇ� �1�'�_�w�}�W�������RF��^�����u�_�u�u�w�p����&�Ə�XF��Z��6���u�u�u�x�!�2��������z��s��!��� �1�'�}�~�}�W���Tސ��\�������!�6�4�4�"�u�^���Y�����X��U����!�;�&�3�2��ԜY���K��X��ʶ�6�;�;�&�3�u����
���OǻN��U���;�0�d�u�9�4�ϩ��ȉ�C"��e�����}��|�u�w�}�WϹ�������FךU���u�u�u��'�����D����F���U���0�0�u�4�0�}�W���J���l�N��Uʥ�'�u�4�u�]�}�W���Y�Ə�XF�N��U���k��8�9��6�W���Y���F���U���
�:�<�_�w�}�W���Y����R/��N��U��6�4�4�:�8�3����0���K��YN�����:�<�
�0�#�/�C�������V�N��U���u�6�4�4�"�}�W���GӅ��G��CF��Y���u�u�u�x�w�(�W���&����P9��T��]��1�"�!�u�~�}�W���Y����r��b �����h�u�:�=�%�`�P���U���F�N��Uʦ�1�9�2�6�!�>����@ӂ��]��GךU���u�u�u���)�������\��U��U���u�u�u�u�w�p����
����\��h�����g�u�:�;�8�m�}���YӃ����R��ʒ�;�%�%�n�]�}�W���K����	l�N��U���e�2�;�'�#�W�W���Y����[	��h�����%�:�;�0�w�2����J���F������u��%��;�$�E���Y�����X��U���u�4�%�0�;�W�W���Y�˺�\	��VN�����;�6�4�4�8�2����0ۯ�F�N����>�4�6�4�6�(�W�������/�N��U���#�:�>�4�4�>��������\��=N��U���x�=�:�
�w��>�������	��R��K��|�u�u�u��(����CӃ��Z��@��[����%�:�;�2�}�%���s���F�P�����8�%�}�u�w�}�W�������w��NN��U���u�x�<�u�>�)��������T��XN�O���_�u�u�u�w�2�ϳ�	��ƹF�N��U���u�u�u�u�w�`�W���	����XJ�N��U���u�x�<�u�$�9�������F�N��1����u�u�u�j�}�3���-����]��~F��Y���x�<�u�&�3�1��������AN��
�����e�_�u�u�w�}�W�������F�S����4� �}�|�w�}�W���Y����F��C
�����
�0�!�'�d�}�������F�N��Uʶ�6�;�;�&�3�}�I�������X�G�U���u�x�u�;�w�)�(�������P��\����!�u�|�u�w�}�W�������G3��D��H���%�;�n�u�w�}�W���Y���F��CN�����2�6�#�6�8�u�NϺ�����OǑN�����2�;�'�!�w�8�E�����ƹ��	�����0��;�:�9�8��Զs���"��V�����4�4�#�9�3�.����Y����R����U���0�<�0�1�;�$�W�����ƹK�r����� �1�'�y�}�3���/����|��=N�����&�}�4�%�2�1�^�������9F������;�
�1�0��0�����Ƹ�VǻN��U���!��9�1�8�3�_���E�Ư�R��V��<��x��!��;�9�������9F�N��Xʘ�&�u�=�u�6�<����Ӊ����^ �����!�u�u�u�4�<��������]�N�U���!��9�1�8�3�_���s���F��V������ �1�g�w�`��������W4��Y
��\ʴ�1�;�!�6�2�8�2���s���V��^�Uʰ�1�%�:�0�$�W�W��Y����G��S��U���<�u�&�7�4�}�Ϫ��״�P
��\N�����y�4�1�4�>�3�ϩ��Ƹ�VF��CךU���!��9�1�"�}�JϽ�����_��X��]���_�0�1���W