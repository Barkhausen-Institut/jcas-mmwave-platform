-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��GZ�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mώ�0����KǶN����g�u� � �#�o�F�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�}�|�g�f�}��������}��X ��U���!� �0�!�w�2��������K��[�����&��&�'�2�W�Zϐ�����_F��D�����&��!�'�6�}��������]l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z��������2��DN�����0�!�<�&�6�)����Y�ƈ�cR�������'�1�3�'�6�}����s����F��^��Uʜ�u�&�1�&�9�8�W����Ư�^��^��U���=��y��{�<�ύ�����HǶN��Dʓ�u�;���]�p�W��?�Ə�9K�N��'���x�_�x�6�4�(�"����ƥ��������1�!�u�0�"�8�W�������`6��B �����u� �u�4�?�/��ԑTӇ��V����U���6�;�u�=�w��C���Y����VF��V�����:�=�'�3�%�)����Y����\��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W��������V��=N�����0�0�&�1�;�:���O�ȭ�_]ǻ��U���0�;�8�'�4�.������ƴF��Y�����!�4�&�4�2�2�������3��d'�����u�����2��������*��C�����0�<�u�'�9�1��������]��NN�����a��1�'�>�}�}�������PNǻN��&���'�6�u�u�#�����Y���A�d�����}�u�u��<�}�W���Y����Z��C
�����n�u�u�6��}�W���Y����Z��C
�����
�0�!�'�c�}�������9F���U���u�u�u�o�>�}��������E��X��Bʱ�"�!�u�|�]�}�W���Y���F�T�� ���!�
�:�<��8����M�ƨ�D��^����u���!�9�.�������G��X	��*���!�'�g�u�8�3���Y����]��F�����1�0�n�_�6�>��������a2��X�����%�m�1�0�w�.�}�������V��S��M�ߊu�u�0�0�>�u�W���Yӧ��`%��pN��U���u�u�o�<�#�:���Y��ƹF�/��8�����u�u�w�}�MϷ�����\�UךU���u���u�w�}�W���Y�����R	��U��d�_�u�u�w��8���<����g2��y1��!���u�u�u�u�m�?�������u'��rUךU���u� �����6���+����g#��h!��<���o�&�'�;�w�`�U���:����F�N��<����u�u�u�w�}�W�������\�*��0���n�u�u�u���4���Y���F�N����2�'�o�u�l�}�W���;����F�N��U���u�o�<�!�0�/�M���B���F��h'�� ���u�u�u�u�w�g��������D��e+��W�ߊu�u�u����%���Y���F������u�h�d�_�w�}�W���+����v*��pN��U���u�;�0�0�w�`�F�ԜY���p4��N��U���u�u�u�u�w�3����Y���l�N��8���u�u�u�u�w�}�W���Y����E��X��Hʍ�f������U�ԜY���~4��N��U���u�u�u�u�w�3����Y���l�N��8��������}�W���Y����T��S��N���u�u�����0���Y���F��^ �����o�u�n�u�w�}�'���<���F�N��U��7�!�#�6�8�}�Jφ�I����V��^�N���u�u���w�}�W���Y���F��^ �����o�u�n�u�w�}�$���4����F�N��U��&�'�;�u�j��6���B���F��r"��4����u�u�u�w�g��������D��c:��;��u�u�u����"���7����`-�N�����u�h�w����<��Y���5��h#��0���u�u�u�u�m�.����Y���`'��UךU���u��
� ��}�W���Y�����^ ��O�����
�w�]�}�W���*����g2��y1��!���u�u�!�<�0�g�W͐�&����v2�=N��U����
���w�}�W���Y����G��PN�UȚ��m�|�_�w�}����s���F��|N��U���u�u�u�u�9�}��������l�N��4���u�u�u�u�w�}�W���Y����_	��T1�����}�l�1�"�#�}�^�ԜY���r%��N��U���u�u�u�;�w�)�(�������P��\����!�u�|�_�w�}�W���,���F�N��U���u�!�
�:�>���������W	��C��\�ߊu�u�u�u�w�}�W���Y�������*���<�
�0�!�%�l�W������]ǻN��U����u�u�u�w�}�MϷ�Yӕ��l
��^�����'�d�u�:�9�2�G��Y���$��b:��U���u�u�o�:�#�.��������V��EF�U���;�:�e�n�w�}�Wϝ�Y���F�N��Oʼ�u�&�1�9�0�>����������Y��E��u�u�u��w�}�W���Y���	F��CN�����2�6�#�6�8�u�@Ϻ�����O��N��Uʅ��u�u�u�w�}�W����ƿ�W9��P�����:�}�b�1� �)�W���s���F��x;��U���u�u�u�u�"�}��������E��X��Bʱ�"�!�u�|�]�}�W���8����}F�N��U���;�u�!�
�;�:��ԜY���p'��n!��U���u�u�u� �w�)�(�������P��]�����:�e�n�u�w�}�4��� ����z(�N����&�1� �:�>�f�W���Yӥ��a?��d-��!���o�:�!�&�3�(����B���F��g#��0���u�u�u�o�>�}��������l��C��Cʱ�"�!�u�|�]�}�W���5����vF�N��U���;�u�!�
�8�4�(��������Y��E��u�u�u����9���Y���	F��N�����2�6�#�6�8�u�W������]ǻN��U�������w�}�MϷ�Y����F
��^�U���u������#���Y�ƣ�GF��S1�����n�u�u�u���1���Y���F��X����� �:�<�n�w�}�Wϋ�=����|1�N��Oʺ�!�&�1� �8�4�L���Y����r2��e ��0����o�:�!�$�9������ƹF�>��!������u�m�2�ϭ�����T��=N��U����d�u�u�w�}�W������G��[���ߊu�u�u��e�}�W���Y�������*���2�6�_�u�w�}�2���4����F�T�����!�
�9�2�4�W�W���Y����F�N��U���u�;�u�!��1����s���F��u\��U���u�u�u�u�9�}��������l�N��6���u�u�u�u�w�}�W���Y����F
��^�U���u������W���Y�ƥ�F��S1�����n�u�u�u���%���Y���F��^ ����� �:�<�n�w�}�Wϝ�4���F�N��Oʼ�u�&�1� �8�4�L���Y����v+��c-��'���u�o�<�u�$�9������ƹF�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U�����u�u�w�}�W������G��[���ߊu�u�u����6���0�������*���2�6�_�u�w�}�$���,����F�T�����!�
�9�2�4�W�W���Y����F�N��U���u�;�u�!��1����s���F��c-��U���u�u�u�u�9�}��������l�N��'�����u�u�w�}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u��	�W���Y���F��^ ����� �:�<�|�]�}��������V��=d��X���%�:�0�e�f�m�F���T�ƭ�F��RN�E���:�u�u�u�m�W�W������W�_�����x���]�}��������r
��X
��Oʦ�1�9�2�6�!�>����Y����G	�N�U��w�s�>� �#�<��������A��d�����_�u�1�%�o��W���
����9F��R �����4�}�u�u�6�<����Y���l�N�� ���0�0�u�k�g�W�W������F��N��U���u�u�u�u�w�}�W���Y���F�NךU��� �:�0�0��<����&����P�	N�����_�u�u� �8�8��������]9��C��*���<�#�h�u��	�?��Y����l��B��K������y�w�}��������X�d��Uʷ�0�u�k�d�]�}�W�������X�s'��6���_�u�u�4�%�4����D����9F������&�9�0�u�i�m�}���Y����[�BךU���4�>�h�u�u��1���?����JǻN�����h�u�y�u�w�0��������A��
P��Y���u�:�8�1�%�:�J���U�����C��U��-�e�e�e�g�m�G���s���C��S�D�ߊu�u�0�
�8�3��������X�d+��8���w�_�u�u�2�����D����r5��d��Uʦ�9�%�!�0�9�`�W͎�-����JǻN����� �!�h�u���U�ԜY�ƹ�V9��C�����!�6�u�k�u��'���<����F�B�����u�k�w��c��}���Ӌ��l�N����u�9�y�u�w�<�J���8������Y��D���_�u�u�u�i�>�5��Y����G	�BךU���u�k�6�y�w�}���� ���F�BךU���6�;�h�u�8�5���^���9F�����u�:�=�'�j�z�P��Y����P��
P�����'�h�r�r�{�}�WϽ�����@��S�R��_�u�u� �#�4����D���JǻN�����u�k�6�6�"�����U�����B��Kʺ�0�y�u�u�4�/��������X��G�����u� �!�<�9�(�W�������9F���Kʶ�y�u�u�%�#�8��������X��G�����u�4�!�'�3�)����GӉ��]JǻN�����9�"�h�u�'�3�}���Y����A ��@N��U���;�_�u�u�6�/����D�ƣ�V�N�����!�h�u�%�9�W�W���	����[�^�E��w�_�u�u�;�0����GӍ��F+��RBךU���4�'�<�&�;�`�W��I��ƹF��R�H���d�y�u�u�4�<�W���^����F�T�� ���0�h�u�d�{�}�WϽ����A��d��Uʶ�7�u�k�r�p�W�W������A��d��Uʶ�6�'�,�;�j�}�F��Y����V�	N��R�ߊu�u�0�!�;�`�W��U�����S�R��_�u�u�0�"�)�������A��d��Uʧ�!�u�k�r�p�W�W���
����^	��S�R��_�u�u�&�5�`�W��U�����TN��U��y�u�u�'�#�1���� ���F�BךU���&�8�h�u�g�q�W�������A
�	N��R�ߊu�u�&�%�j�}�G���Y���9��<��N�