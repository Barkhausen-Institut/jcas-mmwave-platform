-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��E)�� ���=�_�x��#�2�MϚ�Ӥ��VǶN�����4�u�'�?�4�g�'���&�޴�9K�s��O��u� � �!�e�l�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����}�|�g�d�w�2�����Ƃ�G��V����� �0�!�u�8�-�������'��<������&�'�0�]�p�9�������z��E������!�'�4�w�3��������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��/����s����[��T�����!�<�&�4�#�<����Y����CF��+��3���=�&�u�:�'�3����YӲ����U��X���3�%�4�0�w�.����V���r ��EN��ʲ�:�%�:�u��}����
ӏ��R��S
��U���0�!�_�x�4�0��������F��C�����=�'�_�x�z�}��������V
��S��0���'�=�&��;�$�\ϵ�����A��^�����_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���Q��NN����u� �0�<�2�s��������W����N��� �0�<�0�y�(����&����R
��=N�����:�>��2�&�<����݇��l��Y��ʐ�%�<��:�'�4�}�������PNǻN��;���=�&�&�u�w�}�MϷ�������P��U���m�o�u�n�w�}����:����V��V��Oʼ�!�2�'�'�9�8�FϪ�Y���F��=N��U���:�%� �u�w�}�W������V��V ��U���:�b�o�u�w�f�WϮ���ƹF��[��U���u�u�u�u�9�.��������F�T*�����u�u�u�o�>�}����=����GN��B�����x�u�:�;�8�m�L���YӅ��G��[�����u�;�&�1�;�:��ԜY�Ư�\��YN��U���o�<�u�:�1�2����B�����R��U���u�u�u�;�$�9�������F��B�����u�u�o�:�#�.��������V��EF�U���;�:�e�u�l�8�ϛ�	����A	��dװ���<�0�!�'�w�	�W���<����A!��B���ߊu�<�;�9�4�9�������\��G�����}��8�=�$�.�FϺ�����O�
N�����&�k�:�=�%�`�P���P���@��V��1�����'�0�w�}����=����GN��B�����x�u�:�;�8�m�W��Q����A������k�e�|�n�]�8��ԶY���w��Y
��ʺ�u�=�6�u�%�(�W�������[��^����'�;�0�!�2�9��������Z��N@ךU����&�u�1�w�8����������(��ʼ�u�=�u��c�z�W�������_�������{�u�!�u�z�}����	����V��DN��ʻ�"�&�u�4�'�8�W���Y�ƥ�	��R�U���u��%�m�"�8����s���K��E��E��u�y�d�u�{�n�W���T�Ƌ�\��R��D���y�f�u�u��q�E���Y���F�(�����u�x��:�'�}�J��Y���F��F�U���u�u�~��w�v�1�ԜY���!��B�I���y�a�u�y�a�}�D���R���M��N�3���_�u�x��>�}����
�ƾ�R��Y	��U���u�4�4�:�3�/����������S
�����-�'�u��y�}�Z�������@F��Y�����u�=�u��>�}����*������C�����3�_�u�0�%�<������ƹ��T��]���!��|�u�5�:����YӀ��/��YN�����8�=�&�$�l����s���F��V�����!�1��u�j�>�����Χ�A	��y��<���:�u��8�?�.���Y����]��X�����;�u�'�6�$�f�}���Tӱ��[����U���<�;�!�u�6�8����	����@F��[N��U���:�0�9�;�y�}�Ϫ�����FǻC����u�:�&�r�w�2�Ϩ��ƻ�_
��X�����2�u��u�2�}�1�������\��
N�� �ߊu�x�3�'�2�>�W���
�Ƹ���T�����!�0�%�4�2�}�Ϫ��Ƹ�V��E�����9�u�;�4�;�3�Y���>����A6��D�����:�u�u�;�g�)�W�������V�	�����0�u�u�x�!�2����<����A6��DךU���x�=�:�
�w���������/������&�&�>�'�"���ԜY���E��\1�����4�;�6�4�6�3����ۯ�F�C�����4�6�:�3�9�>����ۯ�F�C�����4�6� �%�#�>����6����l�N����>�4�6�:�1�8������ƹF��F�����&�-�u�;�>�$� ���W����Z��V��]���|�u�u�u�0�3�������9F�N��U���8�:�3�0��<���Y����p	��g�����y�u�u�u�w�}�Z����ƥ�G��EN�����d�!�u�m�m�}�}���Y���X#��E�����u�u�u�k��`����)����@K��E��;���|�u�x�<�w�?�������U��Rd��U���%�'�u�4�w�W�W���Y�Ə�XF�N��U���k��>�u�w�}�W���Y���K��YN�����:�<�_�u�w�}�W�������F�S����4�;�:�!�3��[���Tӏ����h�����0�!�'�d�w�2����I���F�N�����4�<��u�i�>��������]J�N��X���;�u�!�
�8�4�}���Y���P%��Q'��U���u�k�6�:�1�3�>��Y���F���U���
�:�<�
�2�)�ǵ�����W��N�����u�|�u�u�w�}�������F�
P��6����y�u�u�w�}�W��Y���@��[�����u�u�u�6�"�-����Y�����S�� ���|�n�u�u�z�}��������T��A�����b�1�"�!�w�t�Wϻ�Ӂ��V��RN������4�0�n�]�}�Z�������v��S
��!���_�u�x�=�8��W���	����P'��R������%�1�0��8����������\@�����0��0�u���}���Y����A��Z��]���u�u�>� ��<����GӍ��^6��D��U���u�;�u�;�2�8�W�������G	�T��A���u�%�'�u�6�}�}���Y�Ə�XF�N��U���y�u�u�u�w�p����
����\��=N��U����%�!�u�i�>����6���K�^ ��&���4�4�!�>�"�����T�ƨ�D��^��U���u�6� �%�#�`�W�������F�C�� ���!�
�:�<��8����M�ƨ�D��^�����;�u��n�