-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��R�����;�{�=�_�z�����CӢ��$��RחXʚ�<�<�4�u�%�7���)����^��=C�1���o�g�u� �"�)�E��s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�}�|�e�l�W��� ����GF��C�����;�!� �0�#�}��������]l�/��U���=�&��&�%�8�}��7����]��~ �����;�&��!�%�<�W�������Z	��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�'�������K��_�����:�0�!�&�:�1�Ϫ�Ӆ��U��N�����9�u�;�u�8�;�Ϸ�Y����`��[�����u�:�4�;�w�<��������G	��_�����0�9�g�u�8�<�����ƪ�]��A�����2�:�!�x�w�2�W���Y����[��F����� �&�u��w�1�ϳ�����V
��R
�����:�&�:�u�?�}��������K��D��U���r�u�:�u�$�}�Ϫ�ӣ��u��_��U���%�;�;�&�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d�����,�<�0�n�w�(�Ϸ��ȿ�W9��P��D��{�9�n�u�"�8����W����A��D�����_�u�&�u�8�6�'�������_
����N���;�<�,��'�2����	������N�����6�_�u�u��0����
���F������u�4�2�u�w�2�O��Y��ƹF��y�����0��4�0�m�4����Ӕ��T���A���h�m�|�_�w�2��ԜY�Ɵ�^��t��U���u�u�u�;�$�9�������F��Z��6���-�u�u�u�w�3��������l�N�����0�3�'�u�w�}�W�������R��N�����3�0�u�u�w�}�W���ӕ��l
��^�����'�g�1�"�#�}�^�ԜY�Ư�\��^ ��U���u�u�u�;�$�9��������G	��Y�����:�e�n�u�w�>�������F�N����!�
�:�<�l�}�WϽ�����z/�N��U��:�!��0����������[��DC����!�u�|�_�w�}�4���-����F�N��U���u�:�3�:�>��_�������V�
�����e�n�u�u�4�2����:���F�N��ʖ�0���'�#�6��������F��@ ��U���_�u�u��2�	�&���Y���\��B�����:�<�
�}��0����
����\��XN�N���u�6�:�3�2�/�W���Y����\��D�����6�#�6�:��}�������]��Y
�����0��8�9�9�f�}������P��RN��9ʺ�u�$��0��0����Y��ƓF�-�����<�;�&�u�#�-�W�������J9��N�����'�4�}�u�8�3���Y����G��X	��*���!�'�>�:�1�4���Y����G	�UװUʦ�2�4�u��2�l�W���Y����@��[�����6�:�}��2�
����Hӂ��]��G��H���!�0�&�k�g�t�}���������R��U���u�u�u�!��2����������R�����d�1�"�!�w�t�M�������@[�I����<�;�9�6�8�;����H�����h�����0�!�'�f�3�*����P���	��R��K��|�_�u�<�9�1��������JT��T�����:�<�
�0�#�/�DϺ�����O�
N�����&�k�e�|�]�}����Ӆ��V ��v�����u�!�
�:�>���������\��XN�U��}�!�0�&�i�m�^�ԜY����R
��t��4���u�u�u�u�8�;����Y���\��E��]���0�&�k�e�~�f�}�������]��t��&���0�u�u�;�2�8�W��Q����c��R��\��� ��0��%�5���s�Ƹ�C�-�����<�
�u�u�$�<����Q����U5��{��Dʱ�"�!�u�|�8�}��������E��X��6����1�=�d�3�*����P���@��V��6����9��u�w�}��������GF��F�����h�}�!�0�$�c�G���B����Z��[N�����'�&��u�m���������\������k�:�=�'�j�z�P���s�ƿ�T�������9��u�u�w�2��������	[�X����}�!�0�&�i�m�^��Yӕ��]��T-�����&��u�o��8�4������F��C����:�=�'�h�p�z�^�ԶYӇ��A��C�����o�&�'�;�l�}����������GN��U���0��,�u�w�}�W���Y�ƿ�T����W���0�n�u�4�#�4��������\ ��t��"���,�u�u�u�w�}�W�������@F��E��N���0�<�_�u�z�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƹK�t�����0�!��4�>�:�4�����ƹK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�x��<�.��������P��C�����'�!�u�;�5�8�����Ə�XW��S�����4�1�!�4�$�8����T�Ƹ�V��XN��ʖ�>�-�1�8�>�s�W��Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d��X���<�&�u�4�'�8����:����R��C��6����u�<�;�;�4�W���Y����_��\N�����{�u�4�>�w�p�W���Y����Z��[N�����:�u�=�u�2�8��������l�t��D���o�u�%�:�2�.�$�������l�U�����u�<�u�<�>�:����Q����_��\G�����u�u�u�6�8�;���Y����U"��d��U���3�'��<�w�}�������F�N�����;�<�;�1�4�2����P������Yd��U���u�u�6�:�1�8����Q���F��X���ߊu�u�u�u�;�8�W���Y�����R��4���-��u�h�p�z�}���Y���V��^�U���u�0�1�9�8�f�W�������U]ǻ��U���6�&�n�_�w�p�9���Y����@ ��������8�9��<�%�������K��[����� �u�=�u�8�;����Y�����^��]���u�0�u��~�;�Ϫ�����A��X ��Uʖ�0�g��o�w�-����
۵��C
��[��\���7�2�;�u�w�4�W�������W��d�����>�-�u�=�9�}�W��������
N�����-�_�u�u�w�p�G��0���/��\��6���h��u�u�w�;�ϗ�����G	������u�u�u�<�w�����!����G��=N��U���u�u��0� ��ݦ�0�����R��4���-��n�u�w�}�Wϻ�
���F�N�����3�0�'�g��t�K���I��ƹF�N�����3�_�u�u�w�}�4���8����F������n�u�u�u�2�9����B���F��t��"���,�6�u�h�4������Դ�9F���U���_�u�;�u�%�>���s�Ư�\��R/��U��6�:�3�0�%���ԶY���z ��g-��U���=�;�"�u�6�}��������F��D��U���4�&�u��9�2����
���Z ��y�����&�z�u�u�2�8����Y���F��^�����:�u�'�4�2�}�%���Y����G��T�����0�!�u�:�w�<�Ϯ����2��DN�����_�u�u�x�#�8�����Ƹ���G�����;�"�0�0�>�}��������F��^�����&�!�8�;�w�<����s���K�=��Y��u�:�3�u�{�e�W���Y���N��G��Yʺ�!� �&�4�2�e�F���O���R�=N��U���3�'�&�_�w�}����
�Ο�^��t���ߊu�u�0�<�]�}�W���Ӕ��Z��R
��]���%�0�9�g�~�)��ԜY���F�^��U���u�h��u�j��W���0���F������3�0�'��;�m�J��Y����K�~'ךU���u�u�u��2�����Q���F��X�����|�_�u�u�w�}�W�������@/��\-������;�d�1� �)�W���E�Ư�\��E��<¾�:�3�'��9�o��������l�N��Uʰ�1�<�n�u�w�}�WϷ�Y����U1��E����h�d�u�=�9�p�W���Y���F������9��}�|�k�}�4���8���]ǻN��U���u��0��;��_���������N�����u�|�i�u��8�$���0�Χ�\��E����1�"�!�u�~�W�W���Y�Ʃ�WF��d��U���u�<�u��2�
�6�������A�������u��u�u�w�}�WϽ�����_��^��I����0��,�e�f�W���Y�����R�����}��0��;�8�Z�������W�S��6����9��}��8�$�������W	��C��\�ߊu�u�u�u�9�}��ԜY���F��������,�6�}�~�z�PϪ����7��N��U���u�6�:�3�%�.�>��Y����p	��v��F��u�u�u�u�w�>����������R�����x�u�:�;�8�l�W������`��f'��6����9�0�x�w�2����I��ƹF�N�����3�_�u�u�w�3�W���s���V��G�����_�u�u�x�w��W���	����@��t��4���u��0��;��^���Yӄ��ZǻN��U���0���}�~�a�W�������V�=N��U���:�u�u�;�f�)�W�������V������u�u�u�6�8�;����0�����R�����}��>� ��8�'�������W�=N��U���;�u�:�%�]�}�W���Y����V��=d��U���u��u�u�'�2��������r�������9��|�u�w�?����Y�����R��<���|�i�u��2����B���F��X��U���d�!�u��:�5����Hӊ��Cl�N��Uʶ�:�3�:���}�JϽ�����_��F������0��'�?�.�^��B���F��Y
�����_�u�u�;�w�/����B���F�?��U���%�:�0�&�4�2����UӅ��V ��[��\���u�7�2�;�w�}�WϽ�����b%�N�U���0��,�g�l�}�W���������N��U���8�=�&�&�f�1��ԜY���F��X������u�h�6�8�;����:�΅�X(��t��%���=�&�|�d�l�}�W�������\	��=N��U���u�'�6�&�l�W�W���Tӷ��F�G�����6�:�3�'�{�>��������l�N�����u�u�u�6�8�;����I�����R����n�u�u�u�1�/�>Ϸ�Y�Ƹ���Z>�����d�9�:�_�w�}�W���:����\7��~G��Hʶ�:�3�'�&��u�]�������c��_��\��n�u�u�u�2�9����B����������n�_�u�;�w�8����ӡ��p	��d��N�ߊu�x��'�#�8�$���Kӓ����RN��U���1�!�u�4�"�1�϶��ƹ�	��NN��ʳ�'�!�#�9�2�}�0���	�ԏ�V ��N��U���8�=�&�&�f�:�������F��X�����e�u�h�6�8�;����P���F��X�����e�u�h�6�8�;����P���F��X�����e�u�h�6�8�;����P���F��X�����e�u�h�6�8�;����P���V��P�����u�0��6��8�L�Զ����g*��