-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��C��&���9�;�{�=�]�p�6�������R��V������<�<�4�w�/����CӶ��V9��OחXʑ�!�o�d��'�8����K����KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��t�E��Y����A��CN�����4�u�;�!�"�8��������R��Yd�U���u�<�=�&��.����s����R��Y��<���'�8�;�&��)����Y����A��^��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��)����@��C�����6�8�:�0�#�4��������G��Q��ʴ�1�'�4�1�$�?�����ƪ�AF��RN�����_�x�3�9�2�}��������F����ʧ� �1�u�=�w�����0�Ƹ�X��^ �����<�u�=�_�z�����:������V�����%�&�0�u�#�)�W���Y����_��\N�����{�u�=�u�9�(�W������Z��E�����&�6�u�=�#�u�^Ϸ�Y����]��D�����u��0�:�#�(�W���ӏ��R��Y	�����&�6�u�=�#�u�^Ϸ�Y����\
��D�����u��<�u�6�>�����ƀ� ��vN�����0�!�!�:�]�p����(ӂ��RHǶd�U���u��a�r�w�.�ϸ�Ӓ����R�����&�7�'�6�8�.��������WF�������u�=�_�x���Oȭ�����U	��C�����1�;�y�4�3�<�����Ƹ�VF��X�����<�6�:�&�9�s�W���
���Z��E�����3�'�8�0�>�:�����ƪ�\��_�����u�-�!�4�$�)���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�<�'�'�w�8��ԜY����Z����*���<�
�d�a�6�1�}���
�ƥ�V��B�����!�{�9�n�w�(�ϩ��Ȝ�T#��V�����4�9�_�0�#�)�W���6����G5��G��ʼ�_�u�0�0�>�u�W�������F�N��U���o�<�!�2�%�/����KӒ��P�
N�\�ߊu�:�!�_�w�}��������F�N��U���&�1�9�2�4�W�W�������p
��ON��U���u�;�&�1�;�:��ԜY�Ư�V��r��U���u�u�u�;�$�9������ƹF��s��<���u�u�u�u�m�4�W���=����GN��d��G���u�:�;�:�g�f�W�������z��N��U���o�<�u�%��)�(�������O�
�����e�n�u�u�4�<�������F�N��U����!�
�}�<�-�X���Hӂ��]��G�U���6�4�4�;��}�W���Y�ƥ�5��s��*���>�%�z�|�f�9� ���Y����9F������9�1�;�u�w�g��������T��=d��Uʶ�4�4� ��w�}�W���Y����|��B�����}��6�d�3�*����P���F��V�� ���u�u�u�u�w�(�W���	����G������1�"�!�u�~�W�W�������e��S!��U���o�:�!�&�3�1����P���WF��G!�����4�%�<�2�]�W��������A��c"��ʐ�%� �%�!�6�-������ƹK��_��*���&�4�!�u�z�+����
����Wlǻ�����6�4�4�1��?�W���Y�Ɵ�P"��V1��]���6�g�x�u�8�3���Y���\��E��]���0�&�k�e�~�f�Wϭ�����P"��V/��&����,�u�u�'�����Qۍ��PI��_�����:�e�u�h��)����Gۉ��V��	I�\��u�&�2�4�w���������F�T�����!�
�}�>�'�r�^������\F��T��]���0�&�k�:�?�/�J���^����F��P ��U���!��1� ��1�W��*����G��F�����|�d�1�"�#�}�^��Yۉ��V��	F�����h�r�r�|�]�}�����Ư�R��X<������u�u�%��)�(���*�����Y��E���h�}�!�0�$�c�������A�d�����4�u��!���������5��s��*����6�d�1� �)�W���C����G��DS����'�h�r�r�~�W�WϪ�	���r��D�����<�u�'�4�w�4����Ӕ��T�N��U���
�:�<�
�2�)���Y����G	�UךU���;�9�6�6�"�����0���	F��t�����!�}��6�e�p�W������]ǻ�����6�6� ��3�/�&���Y�ƍ�p��V
������6�g�x�w�2����I��ƹ��Y�����'�8�:�;�2�.�W�������R��CF�����u�:�;�:�g�f�Wϭ�����P'��E�����0�&�u�u�4�<����&�Χ�C�
�����e�n�u�&�0�<�W���-����]��D'��U���6�4�6�1��u�$���Hӂ��]��G�Uʦ�2�4�u����������\��T-�����
�}��6�f�9� ���Y����9F��^	��ʶ�4�4�4�<��9����Y����_	��T1�����}�u�:�;�8�m�W��Q����A�^��N���&�2�4�u��)�!�������WF���*���<�
�0�!�%�n��������\������k�e�|�_�5�:��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�U���u�1�0�&�6�9�$�������Al�C��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�.�Ϛ�)������t�� ���6�4�4�;��p��������9F�d��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}��������G	��d������<�u�u�8�u�$���K����T��E�����u�x�#�:�<�8�2���
����W��=�����!�'�_�u�w�p����&�Ƨ�F��V��R��u�u�x�#�8�6�ϝ�ӵ��C
��[�����u�x�=�:��}�6���=����]7��~GךU���x�=�:�
�w���������/�N��Xǣ�:�>�4�6�w���������/�N��Xǣ�:�>�4�6�4�(�"����Ư�P)��v
������_�u�u�"�)��������]��NN�����$��%�m�3�8�Wǌ�5���F�P�����8�%�}�u�w�}�Wϵ�����P�	N��R���x�u�;�u�#�����Y���AǻN��U���!�8�%�}�w�}�W���:���F�N��H���4�%�0�9�e�q�W���Y���Z�D�����6�u�u�u�w�>�5���Y���F�������}�|�u�w�}�Z����ƿ�W9��P�����:�}�b�1� �)�W���Y���F��tN��U���u�u�h�u��)�>���Q���F�C����&�1�9�2�4�+����Q����\��XN����u�u�u��w�}�W���Y���P"��V/��&���}�|�u�u�z�2�ϭ�����Z��R����u�:�;�:�g�W�W���Y�Ư�P)��b �����k�6�6� ��9����0����K��B�����:�<�
�0�#�/�E�������V�=N�����0�0�4�0��3��������@]ǑN�����0�&�_�u�8�}�W���IӒ����TA�X���0�0�4�0�]�}�W�������VF��G*��AҔ�1�'��1�%�W�W���T����X9��\=�����!�r�r�u�w�p��������_��V�����g�_�u�u�z�5����Y����P"��V'��6�_�u�u�x�?�2�(���:Ӆ��G��f'��\���u�x�#�:�<�<����=����W��U?��\���u�x�#�:�<�<��������@��T/�� ���1�'���]�}�W�������V��C������%�&�a��9����-��ƹF�	�����u�4�u�_�w�}�W���*����R��
P��E���u�x�<�u�$�9�������V�N��Uʥ�'�u�4�u�]�}�W���Y����F�N��U���8�9��<�%�W���Y�������*���<�_�u�u�w�}�6���Y���F�	N�����;���y�w�}�W������G��X	��*���!�'�a�u�8�3���s���F�T-��U���u�u�u�k�4�<����0ۯ�F�N�U���u�!�
�:�>���������W	��C��\���u�u�u�6�w�}�W���Y�����C�������y�u�z�}��������T��A�����b�1�"�!�w�t�W���Y����r��C;�����h�u���#�9����Q���K�X�����9�2�6�#�4�2�_������\F��=d�����2�;�'�!�w�8�6�����ƓF��R��1���o�u�%�:�2�.�$��������N�����u�u�<�u�>�4�����Ο�^��t�����=�;�u�u�w�>��������z"��R�����4�1��7�l�}�W�������r��B�����h�6�4�4�3����Y����]��QUךU���u�'�6�&�l�W�W��=������
��ʣ�9�1�&�2�6�}�ϳ�����[��^�����1�9�,�}�~�2�W���s���#��s��M���0�&�u��#���������	l�G������8�9��<�%�}�������F�^�����2�0�2�}�6�-����K����[��N��Uʶ�4�4�4�<��9����P���P"��V8�����n�u�u�u�4�<��������`��G��Hʶ�4�4�4�<��9����P���F��SN��N���0�1�%�:�2�.�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�CךU���� �1�'�{�;�ϻ��Ƣ�^�������3�6�0�!�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�CךU��� �0�u��c�z�W���������'�����u�4�4�u��4�W�������R
�������=�u�4�4�w�p�W���Ӓ��G��d�����>�1�8�<�y�}��������Z��^��ʠ�0�u�:�u�!�3�Qϱ����F��Z��U���6�0�3�6�2�)������������ʥ�%�9�;�u�>�;����ӏ��P	��R�����x�u�:�u�'�)����s���9F�N�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x�w�<�Ϫ�Ӵ��]��DN��U���=�u�0�!�#�}�����ɟ�QF��gI�����!�8�;�u�"�-����Y���g��v
��ʺ�!� �u�:�$�)�W���Y����W��^ �����u�4�0�!�2�<����=����V��N�U���!�0�3�'�#�/����Ӣ��F��SN�����=�!�;�-�w�2����
����WF��B ��ʑ��u��&�6�8��������9F��E�������!�1�2�.�[Ͻ�����W��D?����'�8�:�;�2�.�[Ͻ�����a	��S��$�ߊu�0�<�_�w�}�Zό�����N��R��4���'�}�|�u�w�p�W�������W�S�����u�f�_�u�w�p�%������O�
N�����}�|�u�u�z�}�������F�/�����d�_�u�u�z���������Z�e�����}�|�u�u�z�}�������F�<�����u�d�_�u�w�p�%������O�
N�� ���'�}�|�u�w�p�W�������Q�S�����0�u�f�_�w�}����Y���������x�u�:�%�w�}�WϽ�����F��E��<���h�6�6� ��9����Qۍ��PI��'�����}��6�g�~�W�W���Y����\4��Y
�����~��6�g�w�`��������F��E��<��u�u�u�6�4�2��������zO�
N������1�'���6���Pޯ�^	������|�_�u�u�w��#�������@7������u�h�6�6�%�0��������zO��N�����9�:�n�u�2�9��������9F�N�����0�1�!�_�w�/����Q����R'��d��1���u��!��3�(�&���UӅ��G��S=��<����!��1�"��}�������F�C��E���h�}�|�"�#�}�W���s���P"��V:�����0��e�u�j�>��������zN��d��Uʶ�4�4�:�:�9�8�&��Y����w��v
�� ���e�n�u�u�z�}�F���D������_N�3�ߊu�u�x�}�~�a�W��Y����W��qd��U���u�f�u�h��t� ���Y�Ɗ�9F�C�]���i�u�e�u�>�5�FϘ�s���U	��~N��U���:�>�%�z�w�2����Y����w��c�� ���'�}�|�i�w���������w
������x�|�_�u�w�}�3���-����]��fF��U��6�4�4�1��?�3���Q����T�~G�U���0�1�9�:�l�}�W��Y���[�G�����e��_�u�w�p�_���E���F��C��U���u�u�x�u�`�}�J���Pӑ��[F��q(ךU���:�u�u�;�����R�Ƹ���TC����_�u�u�u��)�#�������zN��R�����4�1��7����B���F��s��!��� �1�'�}�~�a�W�������`����ǜ�n�u�u�0�3�1���YӃ����T��N�ߊu�0�� �3�/�M���������N��U���6�d�2�;�%�)�}���Yӡ�� ��RTךU���3��e�2�9�/��ԶY���K��_��*���$��%�:�9�8�W�������9F�N��X���:�
�u��'�����J���F������u�9�u�4�'�8��ԜY���K��X��ʶ�4�4�;�6�6�<��������/�N��U���#�:�>�4�4�<����Y����R)��~F�����u�u�x�=�8��W���6����F����3���� �1�'���}���Y���E��\1�����;�;�&�1�4�>��������zN��=N��U���:�;�0�d�w�3��������v��D�� ���'�}��|�w�}�W�������Z��V�����u�u�u�u��-�3��� ��� O�C�����;�0�0�u�6�:�W������F��N��U���%�'�u�4�w�W�W���Y���p
��N��U���u�k��8�;�����Y���F�C����&�1�9�2�4�}�W���Y����w��~ ��U���h�u��!�������΅�F�C�����!�
�:�<��8����M�ƨ�D��^��U���u�u�u�6�6�<����Y�����C�����|�u�u�u�w�}�Zϱ�ӕ��l
��^�����'�f�u�:�9�2�G�ԜY���F�T/�����&�1�u�k�4�>��������zN��N��U���<�u�&�1�;�:��������_��X����_�u�u�u�w�}�6�������V�	N�����8�:�;�0�$�u�^��T�ƣ�GF��S1�����#�6�:�}�n�9� ���Y��ƓF�N����>�0��%�$�����Ӵ��]��d��U���x�#�:�>�6�6�������� l�N��Xǣ�:�>�4��<�����:��ƹF�C�����
�u��!��}�3���-����]��fF�����u�u�x�=�8��W���������C�����|�u�u�u�z�+����Ӆ��|��Y��ʶ�6�'�8�:�9�8����P���F������u��� �"�8�W���-����]��D?��\���u�u�� �3�/�Mϻ�����D	��+��1���:�;�0�u���}���Y���T��E�����}�u�u�u�w�}��������JF�]��U���<�u�<�!�0�/��������\F��S�����u�u�u�:�#�0����Y���F�-��U���u�u�u�h�w�<�������F�N��U���u�;�u�!��2��ԜY���F�T*�����u�u�u�k�4�<��������A7��B��U���<�u�&�1�;�:��������Q��X����_�u�u�u�w�}�3���6���F�	N����� ���y�w�}�W���T�ƣ�GF��S1�����#�6�:�}�g�9� ���Y��ƹF�N��U���� � �0�w�`�W���-����]��D?��\���u�x�u�;�w�)�(�������P��\����!�u�|�u�w�}�W�������G3��D��H�����:��"�9����0����K��B�����:�<�
�0�#�/�E�������V�=N��U���u�0�0�4�2��ܮ�	��ƓF�p�����o�u�u�<�w�r�GϹ�����VlǻN��U���=�:�
�u�&���������a	��S�����u�u�x�=�8��W���	����R�=N��U���x�=�:�
�w�1�W���	����Xl�N��Xǣ�:�>�4�6�6�<�Ͻ�����a	��S��]���u�u�u�x�!�2��������|��T*�������_�u�w�}�Z�������P'��B�� ���u���:��(����0ۯ�F�N����>�4�6�6�9�3��������a	��S��<�_�u�u�u�8�3���Y����G��X��0���&�� �1�%�u�#���Y���F��R �����4�u�_�u�w�}�W���)����V
��S�G���x�u�;�u�9�8��������F��]��H��u�u�u�u�'�/�W���Y���F�N��6���u�u�u�u�w�c�$�������F�N��U���u�x�<�u�$�9�������F�N��1����u�u�u�j�}�3���-����]��~F��Y���x�u�;�u�#�����&����\� N�����u�|�u�u�w�}�WϽ�����GF�N��U���!��!�}�~�}�W���Y���	����*���<�
�0�!�%�n�W������l�N��U���6�6�;�;�$�9�W�������a	��S��<�y�u�u�x�>�}��������l��C��G���:�;�:�e�]�}�W���Y�Ư�P)��b �����k�6�6�'�:�2����
�΅�]�N��ʦ�1�9�2�6�!�>����@ӂ��]��GװU���u�x�#�:�<�8�2���
����]��<�����a�u�u�u�z�+����Ӎ��C��[��G���u�u�x�#�8�6�ϝ�ӵ��C
��[ךU���u�x�=�:��}�3���0�Ư�R��X<�������_�u�w�}�Z�������P"��V!��U���!��!�}�~�}�W���Tސ��\����:���;�&�1�6�4�/��������bN��=N��U���x�=�:�
�w��>�������P'��X<�����&�}�|�u�w�}�%���������^�����{�$��%�8�3����+���F�N�����'�6�8�%��}�W���Y����c��s����u�|�u�x�>�}��������R��\����o�u�_�u�w�}�W���Ӌ��NǻN��U���u�9�u�u�w�}�W��Y����_��\B��U���u�u�u�x�w�3�W���&����Pl�N��U���6�4�4�;�w�}�W�������g	��B �����|�u�u�x�>�}��������l��C��A���:�;�:�e�]�}�W���Y�Ư�R��B��U���k�6�4�4�"��>��Y���F�N��ʦ�1�9�2�6�!�>����Iӂ��]��GךU���u�u�u�������Y���P'��X<�����&�}�|�u�w�p�W���Y����_	��T1�����}�l�1�"�#�}�^���Y���F��v�����&�1�h�u����������@7��G�X��� �u�!�
�8�4�(������
F��@ ��U���_�u�u�;�w�8����ӡ����RUװUʰ�1�2�;�'�#�}��������@]Ǒ=N��Xʑ�9�,�!�0�3�)�W����ƿ�T�������=�!�0�%�'�1��������	��C��U���u�$��%�o�2����
���w��a�����o�u�%�:�2�.�$�������l�U�����u�<�u�<�>�:����Q����_��\G�����u�u�u�6�6�<����+����V�S��1����9�1�1��?�F��Y���K�z��U���u�4�4�#�;�9��������TF��D��U���u�6�4�4�6�4�%������[��s��#���1�:�;�}�~�W�W���Y����R0��^
�� ���g�u�h�6�6�<����+����W�V �����6�0�0��#�W�W����ƥ�l�R �����0�&�_�u�z�}�����ƨ�G��V��U���7�6�u�;�#�8�F�������W	��^ ����4�<�;�1� �)�W���Y����9F��s��#���1� �u�h�4�<��������]�Uװ�����_