-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��g�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mώ�0����KǶN����g�u� � �#�o�F�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�}�|�g�f�}��������}��X ��U���!� �0�!�w�2��������K��[�����&��&�'�2�W�Zϐ�����_F��D�����&��!�'�6�}��������]l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z���������R��P�����3�'�!�0��/����Y����Z
��E@חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�1���� ӯ��vJ��X�����&�u���$�9��������H��[UךU���u���;�:�/����݇��l��V�����>���'�;�8�W���s���"��VN�����:�u�=�u�o�?�ϱ�����	��C��1���m�&�u�!�'�}��������Z��E��U¼�!�2�'�'�9�8�K����ƿ�W9��P�����:�}�b�1� �)�W���s���F��C�����3�'�!�0�f�}����������C��1���m�&�u�!�'�}����=����GF�������<�!�2�'�%�3���PӉ��@��[�����6�:�}�b�3�*����P��ƹK�s��U���0�3�'�!�2�n�W���Y������\N��U���}�z�y�d�w�3�[��Y����l�C��U���%�!�4�4�#�4�W�������]��R�����u�k�u�3�$�9��������G	��^�����:�e�n�_�w�p��������]��^
��[���3�,� �6�6�:�W���
�Ƶ�FF��A��ʠ�1�!�u�=�w�2�ϳ�	���F��+�����9�9�:�u�8�0����s�Ư�]��Y��6����1�=�u�w�3����Y���]ǻC�1���u�,�0�3�%�)�Ͻ��ƨ�G��XN��ʲ�:�%�{�u�#�-�W�������A9�������,�}�;�0�2�}����Y���\ ��C
�����
�0�!�'�<�2��������W	��C��\�ߠu�x�u�4�6�)�����Ƹ�VF��gZ����1�u�:�!�8�W�W�������|��S��U���&�1�9�2�4�+����Q�ƨ�D��^����x�u� �6�>�3�W���Y����Z��C�����'�6�u�3�#�8�3���Aԕƹ ��T��ʒ�!�&�a��"�>�_�������Q	��R��U��� �;�&�'�9�f�Wϸ�����]F��C*��Aҗ�0�&�>�<�$�g�������A��E �����0�n�u�3�9�)��������^��Z��]���'�!�u�:�;�<�^Ϭ�����|��S��N���3�;�!�:�w�.��������V��^ �����u�0� �;�5�2����s�ƪ�]��X �����1�'�'�0�2�<�_�������V��y�����0��4�0�m�4�����ƾ�G�������n�u�3�;�#�2�W���)����p	�������3�u�;�0�2�t�����ƥ�G��EUװ����6�4�0��:��������l��V�����:�,��2�&�<����ӏ��9F�N�����:�u�:�u�2�)�����ƫ�]��T��ʡ�0���m�$�}��������t��D�&���6�}��'�#�}��������V��YN�����u�&�u�7�0�3�W����Ƨ�Z�������u�u�'�!�%�}�3���:����F�R�����u�u�0� �9��6���=����F�R ����u�0�1��#�.�C׍�����9l�C�� ���<�;�3�'�$�)��������V��^�����=�u��a�p�W�W�������!��s��M���2�}��'�#�}��������V��YN�����'�<�_�u�2�4�}���Y����u��CN���ߊu�u�u�0�"�3�F�ԜY�Ʃ�@ǻN��U��� �;�g�_�w�}�������V��p�����0�&�_�w�p�W������� �������u�=�u�0�2�4�ϱ�Y����w5��I��Uʳ�;�!�:�u�2�����	������E��U���9�4�|�'�#�/�W���������N�����u�u�<�u��/�Ϫ����F�E�����%�:�0�!��m�G��H����K��
/�����u�9�0�u�w�}�����ƃ�^	��h��W��e�e�w�n�z�}�J���R����9F���U���_�u�;�u�2�����	����lǻC�3���!�:�u�:�w�8����Y����T��E��U���!�0���o�.�Wϸ�����]F��r��]���8�0�o�<�#�:����������[��U���u�7�2�;�w�}�����Ƨ�F��EN����h�e�_�u�9�}������ƹK�q�����u�:�u�0�#�3�W���Y����JF��E��ʴ����:�'�.����Ӓ��Vl�Q�����u�0��1�%�/�����Χ�F��V��Y���8�:�3�0��<�������V�E�����;�0�0�u�$�}�WϨ�����VF��S�����u�;�0�0�l�}���������\ ��%���0�h�u�=�9�}�W���8����w
��S��N���u�0�&�3�<�(�'�������G��=N��U���1�0��,�m�}�L���YӃ��Z ��y�����&�a�!�0�]�}�W�������_�
N����u�9�0�u�z�����
���9F�N������,�o�u�l�}�Wϻ�ӏ��9F�������0��'�?�.�J�����ƹF�/�����,�o�u�1�2����s���V��^�U���'�!�'�u�3�8�3���s�Ʃ�WF��C/�����0��9�,�]�}�Z�������\��X�����;�u�=�u�?�.�W���Ӆ��Z��R �����3�;�!�:�w�8�'���������Z-����<�!�2�'�w�8��������V��Dd�����;�u�u�<�w�.��������\�������u�u�'�!�%�}�9�������F�R�����u�u�0� �9�6��������9F���U���_�u�;�u�2���������9l��SN�����0�7�1�u�<��'�������9