-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��S�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������Kl�*�����b��2�&�w�m�B��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���u�6�u�e�b���������R��Y��<���'�8�;�&��/������ƴF��[N�����u�0�0�#�3�p�W�������/��C�����u�;�0�;�;���������9K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x�x�w�(����C���g�������;�u�;�!�9�4����=������DN�����y�!�u�1�w�2�������J��EN�X���$��'�=�$�}������ƴl�>�����0��9�,�]�p�W��*����VǶN��Aʆ��u�g�x�w�}�W���C����K�_�&���u�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��Ɠ_��V�����n�u� �0�>�8�Y���&����P9��Z����u� �0�<�2�s��������WH��[UךU���u�:�>��0�,��������_
��=������%�1�0��8�W���YӁ��V��d��Uʾ� ��4�0�w�}�����ƾ�]��N��U���h�a�|�_�w�2��ԜY�Ə�XF�N����!�
�:�<�l�}�WϽ�����\��YN�����4�!�>� ��<���Y����G	�UךU����!� �u�w�(�W���&����P9��T��]��1�"�!�u�~�t�}���Y����W��c��N�ߠ4�6�<�0�#�/�W���Y����B��S�����<�_�u�x�!�2��������Gl�C�����&�2�;�_�w�.����Y����@��V	�� ���u�%��!��u����)����@I��_�����:�e�u�h��)����Gۉ��V��	I�\��u�&�2�4�w�����*����|��N�����4�!�d�1� �)�W���C����G��DS����'�h�r�r�~�W�������t��d�����_�u�3�>�"�����D�ƫ�]��CךU����!� �u�j�>����
���9F��Y
�����4�0��;��>����s����V��G����u�<�u��:�5����KӁ��V��RdךU���x�=�:�
�w�,�3���A����AF��G*��AҔ�1�'�d�u�w�p��������`��E��U��_�u�u�x�?�2�(���8�Ư�]��DF����u�x�=�:��}�4Ͻ�����W�N��Xǣ�:�>�4�6�w�����s���K��X��ʶ�6� � � �2�}����Y����B��GZ�����-�o�0�!�#�}����<����CR��S
��U��_�u�u�w�8����Y����l�N��Uʾ� �!�4�!�j�}�G���Y����]F��C
�����u�h�r�r�w�}�WϮ��ơ�CF�N��U����>�u�u�w�}�W���:���F�N��X���;�u�!�
�8�4�}���Y���P'��N��U���u�k�6�;�"�.�G��Y����]F��C
�����
�0�!�'�c�}�������F�N�����u�u�u�u�w�c�������J�C�����!�
�:�<��8����M�ƨ�D��^��U���u�u�6�u�w�}�W���Y����|��B�U���x�u� �u�#�����&����\� N�����u�|�u�u�w�}��������@��
P�����n�u�u�u�z�}��������T��A�����l�1�"�!�w�t�}����ƫ�]��C�����%��&�n�]�}����	����V\ǻ������4�0�h�w�8�������!��q�����2�o�u�u�1�/�>Ϸ�Y�Ƹ�W��R �����_�u�u�u�z�5����Y����@��v
��ʐ�%�&�a��3�/�E���Y�����X��U���7�'�6�u�g�W�W���Y�˺�\	��VN��7ʶ�;� �&�g��W�W���Y�˺�\	��VN��U���%�!�}��|�t�W���Y����[	��h��%ʶ�<�&��4�2�(�_���Y���K��_��*�����!�;�$�9����s���F��G*��AҔ�1�'�g�u�9�4�ϩ��ȉ�C"��V�����}��|�u�w�}�WϹ�������FךU���u�u�u��5�/����G����F�N��Uʦ�1�9�2�6�m�}�G�ԜY���F��E�����_�u�u�u�w�}����Y���F�	N�����u�u�u�u�w�}�W��Y���@��[�����u�u�u�u�4��W���Y���X��~ ������|�u�u�w�}�ZϷ�Yӕ��l
��^�����'�a�u�:�9�2�G�ԜY���F�T-��U���u�u�u�k�4�3����Kٯ�J�N��Xʼ�u�&�1�9�0�>����������Y��E�ߊu�u�u�u�w��W���Y���[�T(�����4�0� �}�~�}�Z����ƿ�W9��P�����:�}�b�1� �)�W���Y���F���:���;�&�1�h�w�-���Y���F�N��X��� �u�!�
�8�4�(������
F��@ ��U���_�u�u�;�w�8����ӡ��u��C=����_�u�u�x�?�2�(�������^��S��0���&�a��1�%�n�W���Tސ��\�������6�u�e�_�w�}�Z�������P'��T(�����4�0� �}�~�}�W������l��tN������4�0� ��t�W���Tސ��\�������%�!�u�u�z�+����Ӆ��|��Y��ʺ�0�_�u�u�&��������� \��Y��ʢ�'�{�$��'�e����Y۴��l�N�����'�6�8�%��}�W���YӍ��Q��T��K��r�u�x�u�9�}��������	[�IךU���u�:�!�8�'�u�W���Y����_�N��U���h�u�9�y�w�}�W���Y���F���U���
�:�<�_�w�}�W���8���F�N��Kʶ�<�&��4�2�(�_���Y���Z�D�����6�#�6�:��j��������9F�N��U���u�u�u�u�w�`�W�������R��B��\���x�u�;�u�#�����&����\� N�����u�|�u�u�w�}����Y���F�
P��:��� �y�u�u�w�}�W���TӉ����h�����0�!�'�a�w�2����I���F�N����� � �0�u�i�2����Y���F�N��U���:�!�&�1�;�:��������_��X����_�u�0�1�0�3����Y����`��V������;�c�%��.�M����Ƨ�F��V��H���0�0�4�0�w�}�0�������G��d��Uʳ�'��<�u�w�2�DϹ�����VlǻN��U���=�:�
�u�&���������v��D�4���'�a�u�u�w�p��������`��E��U��_�u�u�u�z�5����Y����P/��B��G���_�u�u�u�z�5����Y����z��C��_���|�u�u�u�z�+����Ӆ��P ��D����� �}�|�u�w�}�Z¨�������x�����1�:�0�_�w�}�W���=����r��E�U���<�,�"�'�y�,�3���A����AF��c"��U���u�u�2�;�%�>����Q���F�N��&���'�6�u�k�p�z�W��Y���@��[����u�e�_�u�w�}�W���Ӌ��NǻN��U���u�9�u�u�w�}�W��Y����F�N��U���u�u�x�u�9�}��������F�N��Uʶ��u�u�u�w�}�IϽ�����T��B��U���u�x�<�u�$�9��������G	��Y�����:�e�_�u�w�}�W���:���F�N��Kʶ�;� �&�g��l�[���Y���Z�D�����6�#�6�:��j��������9F�N��U����u�u�u�w�}�J���?����`��R!��]���u�x�u� �w�)�(�������P��Z����!�u�|�u�w�}�W�������G3��D��H���%�;�n�u�w�}�W���Y���	����*���<�
�0�!�%�o�W������lǻN�����0�0�4�0��3����*����lǻN�����6�;��4�2�W�W����ƅ�Z���Dʲ�;�'�!�_�w�}�W������l��F�����1�0�u�$��-�O�������F�N����>�4�>� �#�<����^���F������u��u��%�)����6���/�N��U���#�:�>�4�4�}�1�������V)��\��^���u�u�u�x�!�2�����Ư�V��S=�����!��_�u�w�}�Z�������P'��B�� ���u�%�;�u�w�}�2���
����W��O[����!�u�:�>��-���8����N��{GךU���u�u�0�0�>�}����s���F�N�� ���4�!�h�u�g�t�W������G��X	��U��r�r�u�u�w�}����Y����l�N��U����>�u�u�w�}�W���:���F�N��U���u�u�u�u�z�4�Wϭ�����ZǻN��U���u��u�u�w�}�W��Y����@��V	�� ����|�u�u�z�}��������T��A�����b�1�"�!�w�t�W���Y�����N��U���u�h�u��%�)����6���/�B��X���;�u�!�
�8�4�(������F��@ ��U���u�u�u�u�w�>�W���Y���F�������4�0� ��t�W���Y����F��C
�����
�0�!�'�c�}�������F�N��Uʶ�6� � � �2�}�Iϱ�����F�N��U���u�u�u�x�8�)��������l��C��G���:�;�:�e�]�}�Wϻ�Ӂ��V��RN�����:�1�!�2�l�W�W���T����X9��r�����1�'��'�.�Cן�����9F�C�����
�u��7�%�>�W��s���K��X��ʶ��6�0�:�3�)�������F�C�����4�6�u��4�3�$�������OǻN��X���:�
�u��4�(����Y�����X��U����!�;�&�3�2��ԜY�Ɖ�C"��V�����c�u�;�<�.�*��������^��S��]���|�u�u�u�0�3�������9F�N��U���7�'�6�u�i�z�P���T�ƥ�F��S1�����o�u�e�_�w�}�W���Ӌ��NǻN��U���9�u�u�u�w�}�J������F�N��U���u�u�x�<�w�.������ƹF�N��4���u�u�u�u�j�}�$�������T��CF�Y���x�<�u�&�3�1��������AN��
�����e�_�u�u�w�}�4���Y���F�	N�����1�!�2��#�l�[���Tӏ����h�����0�!�'�a�w�2����I���F�N��U���u�u�u�u�i�>�������F�N��U���u� �u�!��2��������R��S�����|�u�u�u�w�>����,����WF�����u�u�u�u�w�}�W��Y����@��[�����6�:�}�l�3�*����P���V��P�����u�0�d��4�<��Զs���WF��{U�