-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B6��V�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mώ�0����KǶN����g�u� � �#�o�F�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�}�|�g�f�}��������}��X ��U���!� �0�!�w�2��������K��[�����&��&�'�2�W�Zϐ�����_F��D�����&��!�'�6�}��������]l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z��������2����������6�:�2����Yӯ��F��V ��:��� �&�4�0�<�-�W�������@��V��U���x�u�=�u�6�-����Y����Z�'�����9�,�!�0�2�<�ϸ��Ɗ�aF��[��ʼ�%�0�0�!�3�p�W���Ӎ��^%��Q>��%���0�>�%�z�w�2����������(��[���_�x�u�u�w�}�W��T���K�C�X���u�u�x�x�]�p�>Ϸ�Y���OF��eN�]���;�<�0�u�z�p�W���T���K�������u�u�u�)�w�p�Z��T���K�C�U���x�x�_�x�w�}�WϢ�Y���K�C�X���x�x�u�u�+�p�W���Y�����~<��U�6�:�&�u�+�p�W���T���F�N��U���x�x�x�x�z�p�Z��T���OF�Kd�U���u�u�u�u�w�}�W���Y���F�N��U���u�_�x�u�w�}�W���T���K�C�X���x�u�u�)�w�!�Z���Y���K��(��U����6�:�&�w�!�Z��Y�ư�K�N��U���x�x�x�x�z�p�Z��T���F�N�����u�u�u�)�w�p�Z��T���K�C�U���u�u�x�x�]�p�&Ϸ�Y���OF��eN�]���;�<�0�u�z�p�Z���Y�ư�K�������u�u�u�u�w�p�Z��T���K�C�U���u�u�x�x�]�p�Z�������]��R��O���u�u�=�u�>�8����������VN�����:�u�3�>�'�}����7����V ��E>���߇x�u�u��3�/����s���F�N��6���_�x�u�u�w�}�'��K���F�V��%��a�x�u�u�w�k�$���Y���9K�N�����;�u�0�4�m�p�W����ƭ���YN�����u�3�6�0�1�>����C����(��t��%���=�&�~�1�2����s��� �������;�8�0�u�1�>��������@\�_�;���:�3�0��6�8�6�������TǶd�U���3�<�<�;�w�2�ϑ�����K�-�����<�;�&�4�2�1����Y����G����ʡ�0�=�2�0�#�4����Y����Y��^ ��X���u�:�;�7�w�����
����R��C��Yʸ�1�}�z��:�2���Y����G��`�����u�u�-�8�;�}����Y����RF��R�����&�u�4�0�]�p�Z���Y����
��S��U���u�:�3�<�>�3��������@��C�����3�0�u�:�#�8��������GǶN�����0�{�u�=�9�.�Ͻ�����]F��C��6����h�d�{�w�5����
ӈ��]����U���6�&�x�u�w�8� ���Y����P	��Q�����{�u��0� �}�����Ư�V��SN�����:�1�{�u��8� �ԑT����@F��R
��ʰ�4�9�u�u�?�;�W���������T�����&�!�0�6�2�;�����ƥ�G	��_חX�����m�&�w��W���Y������R��U���=�3�'�!�8�1�������\��^�����"�9�_�x�w�6��������]��Y
�����%�<�u�=�w�/����	����F�������:�1�y�!�2�9��ԑT����]F��X����� �<�2�!�2�1����7����V ��N��ʢ�0�u��0� �`�F���
ӓ��WF��Ed�U���=�u�:�3�>�4����s��ƴF�T-�����_�x�u�u�g�m�W�����ƴF�I�D���u�u�;�<�2�u�>�ԑT���V��N��<ʶ�:�&�u��~�p�W���^����[�������}��_�x�w�}�F��Y�Ɲ�Z��Y��$���x�_�x�8� �+�W�������R
��R��U���u�4�0�_�z�}�$���D����N��B�����h�|�x�u�<�(�4���)����R��
N�]���:�3�<�<�9�.�������F��G�����0�4�u�u�g�����:����J��Dd����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W��������V��=N�����0�0�&�1�;�:���O�ȭ�_]ǻ��U���0�;�8�'�4�.�������F��@��[�����'�9�2�s���s����G��F>�����9�<�2�0�8�}��������Z�N�����u�u�u�u�w�}�W�������AF��Y	��Gʡ�u�c�o�u�a�W�W���7����V ��E>�����u�;�0�0�w�<����Y���F��_��N���%�'�}�u�w�����:���F�N����!�
�:�<�l�}�Wύ�����_��N��U��<�u�!�
�8�4�L���YӅ��@��N��U���u�o�<�u�#�����B�����R�����u�u�u�o�>�}��������E��X��Bʱ�"�!�u�|�]�}�W�������F�N��U���;�&�1�9�0�>�}���YӅ��G��N��U���u�u�;�&�3�1��������AN��
�����e�n�u�u�4�<����Y���F������9�2�6�#�4�2�_������\F��d��Uʶ�4�4�;�u�w�}�W���ƿ�W9��P�����:�}�b�1� �)�W���s���P"��V'��U���u�u�o�<�w�)�(�������P��_����!�u�|�_�w�}�3���0���F�N����!�
�:�<��8����H�ƨ�D��^����u��!��b�}�W���Y�ƥ���h�����0�!�'�d�w�2����I��ƹF��s��<��u�u�u�u�w�3��������l��C��D���:�;�:�e�l�}�WϽ�����F�N��U���;�&�1�9�0�>����������Y��E��u�u�6�4�6�3�W���Y�����D�����6�#�6�:��j��������l�N�����;�u�u�u�w�g��������T��A�����b�1�"�!�w�t�}���Y����R/��N��U���o�<�u�!��2��������W��S�����|�_�u�u��)�>��Y���F��^ �����:�<�
�0�#�/�F�������V�=N��U���!��d�u�w�}�W���ӕ��l
��^�����'�d�u�:�9�2�G��Y����w��~ �U���u�u�u�;�$�9��������G	��Y�����:�e�n�u�w�>�������F�T��ʦ�1�9�2�6�!�>����Nӂ��]��G�U���6�4�4�;�b�}�W���Cӏ��@��[�����6�:�}�b�3�*����P���F��V������u�u�u�w�3��������lǻN��1����!�u�u�w�}�W���Y����_	��T1�����}�e�1�"�#�}�^�ԜY�Ư�R��B�U���u�o�:�!�$�9��������G	��^�����:�e�n�u�w�>�������F�T�� ���!�
�:�<��8����J�ƨ�D��^����u��!��#�}�W���Y�ƣ�GF��S1�����#�6�:�}�g�9� ���Y����F�T*�����a�u�u�u�m�2�ϭ�����Z��R����u�:�;�:�g�f�W�������|��N��U���u� �u�!��2��������U��S�����|�_�u�u��)�8���Y���F��X�����9�2�6�#�4�2�_������\F��d��Uʶ�4�4� �b�w�}�W������G��X	��*���!�'�f�u�8�3���B�����C�����u�u�u�u�"�}��������E��X��Eʱ�"�!�u�|�]�}�W�������
F�N��Oʺ�!�&�1�9�0�>����������Y��E��u�u�6�4�6�(�F���Y���	����*���<�
�0�!�%�n�W������]ǻN��1����!�d�u�w�}�W���Y����_	��T1�����}�e�1�"�#�}�^�ԜY�Ư�R��B�U���u�o�:�!�$�9��������G	��^�����:�e�n�u�w�>��������F�T�� ���!�
�:�<��8����J�ƨ�D��^����u��!��#�i�W���Y�ƣ�GF��S1�����#�6�:�}�g�9� ���Y����F�T*�����d�u�u�u�m�2�ϭ�����Z��R����u�:�;�:�g�f�W�������e��S!��U���o�:�!�&�3�1����s�����V
�����%�!�u�o�8�)��������O��=��U���4�4�9�9�>�:����B����A��C�� �����:�u�&�<��������_��GN�����x�#�:�>�$�:����s���E��\1�����_�_�u�:�$�<�ϵ�����@��N����2�'�o�u��>�E�ԶYӕ��]��T<�����!�u�u�o�$�9�������V�=N�����9�6�0�0��$�W���Cӕ��l
��^��H��r�_�u�<�9�1��������]�T�����;�1�m�1� �)�W���C����G��DS�E���_�u�&�2�6�}�#�������F�N�����;�o�u�4�$�f�Wϭ�����P2��P�����u�o�7�:�2�3�M�������9F��^	��ʶ�:�2�0�3�2�o�Mϼ�����\�Q���ߊu�<�;�9�4�3�������\��X�����h�3�9�0�]�}�Z�����ƹ��Y�����3�:��u�w�g�4���-����l��y�����&�d�1�"�#�}�^��Yۉ��V��	F�����h�r�r�|�]�}����Ӆ��V ��v��U���u�!�
�:�>���������\��XN�U��}�!�0�&�i�m�^�ԶY���w��=N�����9�6�4�4�9�}�W���Y����G"��V1��D���:�;�:�e�w�`�_������	��R��K��|�n�_�u�>�3�Ͻ�����t��G��U��� ��!�
������
�����Y��E���h�}�!�0�$�c�������A�dךU���;�9�6�4�6�2�������5��s��*����8�=�&�$�l��������\������k�:�=�'�j�z�P���s����Z��[N�����'�8�:�;�w�}��������l��d��Dʱ�"�!�u�|�m�}�������\��E��R��|�_�x�u�>�3�Ͻ�����\��B ��U��� �%�!�4�6�)����T�ƨ�D��^��O���:�=�'�h��)����G���]ǑN�����u��!��#�8����Y�ƃ�G��s��*���`�1�"�!�w�t�M�������@[�X����r�r�|�_�w�p�W���
�ƨ�_����U����8�9��<�%����
����\��V ����� ��9�,�w�}�MϷ�����\�U��Xʰ�!�4��u�8�}����Y������X�����:�u�;�>�>���������F��Y������'�=�&��1����Y����T��S�����4�0�:�3�<�(�4���)����R��E��N���6�;�!�;�w���������_��N�����'�o�u�0��9��������JN��B�����y��8�:�1�8�'�����ƹ��D��ʾ�1��7�0�6�}�W������V�
N����:�&�4�!�<�2����=����F������u�h�`�_�w�p�W�������JF��C�����=�u�0�4�w�3�$���������\ךU���&�4�!�>�6�<����)����	F��C����u�>�;� ��1��������[��s�����>�1�0��2�����Y���F�N��U���u�u�u�u�w�}�W���Y���F�\/��&���0�4�u�u��(��������T��=N�����9�6�4�4�6�4�3������	F��S1�����#�6�:�}��/����=����W��X����u�h�}�!�2�.�I��P���@��V��1����9�1�1�2����
����\��h�����>�1�0��2���������\F��T��]���0�&�k�e�~�W�Wϭ�����P"��V8�����:��u�u�w�)�(�������A��d�����4�u��!��1��������\��C
�����u�h�r�r�]�}����Ӆ��G��[����� �&�o�&�3�1����C���]ǑN����� �0�>�0�w�}�������R��^��ʾ�0�u�3�6�9�?�������F�T�����9�<�u�!�"��}�������F��Z����� �o�<�!�0�/�}�������F��Z����� �u�3�6�9�?���������Y�����c�_�7�2�9�W�W��Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=N��Xʖ�0�!�u�;�2�<�������� �������u�=�u�4�6�;����������C��G���9�6�_�u�z�9����W���F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠu��0�!��<����C����A	��D�����0�9�|�u�5�:����Yӏ��A��Y	������8�9��<�}����Y�����P	��3���h�;�!�6�8�:����s���V��^�Uʰ�1�%�:�0�$�W�Wϝ�����]��R\�����'�6�&�}�6�-����K��ƹ��^ ךU���3�'�&�;��9�Ǎ�����_��N���ߊu�u�u��0�1�1��������P	��3��u�u�u�6�8�:�������F��X	�����0�n�u�u�w�>��������F�
N�����0�3�0�g�/�/��������w��=N��U���u�3�_�u�9�}����
��Ɠ9F�N�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x��8��������\��Y	�����<�_�u�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���2��R��ʶ�0�3�6�0�#�}��������V��[��ʡ�0��>�-�3�0�������A��Q�����x�!�0�u�8�)�ϝ�����\��Y@ךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z¨�����#��t��&���9�;�_�u�z�5����Y����U5��L�D�ߊu�x�=�:��}�4���-����\��=N��X���:�
�u��2�	�&���	��ƹK��_��*����0���w�-����<����V ��Z�����u�;�<�,� �/�Y���:����R��^ ��]���|�u�u�2�9�/�ϳ�	��ƹF������&�&�u�u�w�`�W�������V�N��U���x�<�u�<�#�:�Ϭ������N�U�ߊu�u�u��:�2����)����[�\ ��6����'�=�&�~�}�ZϷ�Yӏ��V�������u�:�a�u�j�e�W���	����^��d��U����8�9��<�}�J�������p
��N��X���;�u�!�
�8�4�}���Y�Ɵ�^��t����u�4�%�0�;�o�[���Tӏ����h���ߊu�u�u��6�1�/���Y����v��[�����u�x�<�u�5�2����Y�����R�����u�k�w�e�u�}�W���Y���Z�D�����6�#�6�:��}�������F�N�����<�u�u�h�w��������F���U���
�:�<�
�2�)���Y����G	�d��U���6�:�3�0�w�}�J���:����VJ�N��X���;�u�!�
�8�4�}���Y�Ư�\��X'��U��u��0���q�W���TӉ��%��Q:�����}��8�=�$�.�FϺ�����OǻN��U���0���u�w�c����U���F�C�����0���%�)����)����@K��S�����|�u�u�u�4�2����:���F��R �U���u�u�x�u�"�}��������GN��B�����x�u�:�;�8�m�}���Y�Ư�\��X?��U��u�%�;�u�w�}�W���TӉ��%��Q:�����}��8�=�$�.�FϺ�����OǻN��U���0���,�w�c��������JO��C����&�1�9�2�4�+����Q�ƨ�D��^���ߊu�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���TӴ��V��O�����u�<�6�<�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�����,� �1�!�4�}�W�������W��X �����y�1�4�&�%�}����Y����Z��CN�����x�u�0�1�g�.��������[��^��ʳ�'�g�>�4�6�<����	�Ư�P
������� �!�3�'�w�p�W���Y����_��
�����u�=�u�'�"�}����Y����[��~<�U���u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W�������V��X �Uʥ�:�0�&��:�1�4���s�Ʈ�T��N�����<�<�2�0�0�u����������Yd��U���6�0�0��.�a�W���
����F�N��U���&�!�r�r�6�9��������A�������u�u�u�6�2�8�4������G	��Y�����}���!��1��������P4��R�� ���9�;�!�|�]�}�W���Y����V��CN�U��n�u�u�u�2�.�Ͻ�����\��	^�����u�u�u�u�4�8�������F��D������&�!�:�9�p�^�ԜY���F��R��0���i�u�d�n�w�}�Wϻ�
���F�N������!�i�u�g�f�W���YӃ����=N��U���u�3�_�u�9�}����
��ƓF��R��3���;� �u�h�9�)��������lǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z���������F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�x�u�2�5�����ƨ�G��Y�����,�u�:�u�6�.����Ӓ��#��d�����'�_�u�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���F��GN��ʼ�%�!�1�!�w�2��������F��[��&���&�8�9�&� �1�W���������B��[���6�4�4�;�g�}�K���=����]V��N�����;�d�u�i�w�����H���P"��V'��G���i�u��!��o�}���=����]N��N�U���!��f�_�w�����Q���[��s��<��_�u��!��u�^���DӅ��G��UךU���!��}�|�w�`��������9F��s��<���|�u�h�6�6�<���YӅ��G��V��U��6�4�4�;�l�}�������F�
N�����;�n�u�6�6�<���P���P"��V'��E�ߊu��!���l�W������z��d�����4�;�d�|�k�}�3���0����9F��s��<���f�u�h�6�6�<���s�Ư�R��YF�\��u��!��f�f�WϽ�����W��R�����4�;�`�_�]�}�Z�������v��Y��&���9�;�u�;�"�����0���K��X��ʶ�4�4�;�6�6�<�ǵ�	����W	��C��\���x�#�:�>�6�>�����Ư�R��X)�� ���u�x�#�:�<�<��������W)�������9�1�'�8�9�}�>�������_��N�����u�:�>��'�3��������TF��c"��U���2�;�'�6�:�-�_���Y����`��N��U���u�u�h�u��>�W���Y���F�C����<�!�2�'�%�3�������\�d��U���>� ��0��/����Y����}��X�����4�0�u�x�w�3�W�������A��RN����m�o�u�_�w�}�������9F�N�����0�9�u�u�w�}�W��Y����_��\B��U���u�u�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u�4�%�0�;�o�W���Y���F��Z��6���-�u�u�u�w�}�W���Y����]F��C
�����_�u�u�u��.����Y���F�S����0��!�u�w�}�W���Y���F���U���
�:�<�_�w�}�W�������U��N��U���k�6�;�7�2�;����Y���F�N��X���;�u�:�9�6�W�W���Y����R/��N��U���u�u�k�6�6�<�ǵ�	����W	��C��\���x�u�;�u�9�(�3���&�Χ�C�
�����e�u�u�u�4�<����Y���F�N��U���!���:�'�q�W���Y���F�N��ʜ�%�!�4�4�#�u�$���V���F��=N��U����!��9�3�3�W���Y���P"��V8�����y�u�u�u�w�}�W���Tӏ����h���ߊu�u�u��#���������C�	N�����4�<���8�-�[���Y���K��B�����:�<�_�u�w�}�3���/����|��N��U��6�4�4�4�>�����P���F�N�U���u�!�
�:�>�W�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d��X����u�<�!�%�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǻC�<���4�!�4�0�<�-�X�������t��GN�����0�!�y�0�4�}����������Z>�����u�x�u�3���������g��\=��Z��� �%�!�u�%�}�����ƾ�F��S@ךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}��������C��d������<�u�u�8�6��������F��Y���ߊu�u�x�=�8��W���?����\��r�����:�%��_�w�}�Z�������X!��B��ʜ�u�u�x�#�8�6�ϝ�ӵ��C
��[�����u�x�=�:��}�4���0�Ư�\��X'��U���x�#�:�>�6�>����Ӆ��V ��v��E�ߊu�u�x�=�8��W�������P"��V:�����&�u�u�x�!�2��������e��S'�����4�4�<���2��ԜY���E��\1�����%�!�6�4�6�2��������l�N������:�%��m�8����Y����#��q�����u���_�w�}�W�������^��d��U���u�>� ��6�8�W���Y�����Z>�����u�u�u�u�z�}��������AF��Y	��Dʡ�u�u�h�a�w�}�W�������\��R�����h�u��8�8�;�������K�^ �����2�'�'�;�2�l����A���l�N��Uʾ�'� ��8�w�}�W���Gӯ�F�N��U���u�u�x�u�9�}�����ƾ�]��N��U���h�e�u�u�w�-�������F�N��6���u�u�u�u�w�c�$��������N��U���x�u�;�u�#�����s���F�T*�����u�u�u�k�4�<��������F�N��X���;�u�;� ��)�(���7����R��_�����:�e�_�u�w�}�W�������Z��S����4�4�<���2���Y����]F��C
�����_�u�u�u�w�����Y���[�T-������u�u�u�w�}�W������\��X(��*�ߊu�u�u�u��8� ���Y���F��X�����}�|�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u�u��!�"�}�W���D�Ư�R��X/��&�����|�u�z�2�ϭ�����Z��R����u�:�;�:�g�W�W���Y����A��)��3���'� �&��]�W�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��N�U���4��9�1�#�}����Y����CǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z���������R��A��ʦ�2�4�u�,�#�8����Y����_��
�����&�0�6�u�%�(�Yϟ�
���K��y*�����4�4�#�9�3�;�����ƥ�C��C����� �%�!�!�w�>����Y����G��T�����x�u�;�7�2�2�W���Y����P��YN�����'�=�&�|�w�4��������@F��D�����:�&�_�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƓF��C�����<�0�_�u�%�>��������p
��OGךU���<�_�u�u�1�/����&����5��G�����|�!�0�_�w�}�W�������G#��
I�U���;�u�u�u�w�>��������@��NN�Uº�=�'�h�r�p�f�W���YӃ��Z ��s��#���1�'�8�;�p�z����s���F�T*�����<��%�9�w�`��������W"��s������4�0�0�6�p�W������F�N��U���u�u�u�u�w�}�W���Y����w��a�����8�;�_�u�w�}�������F��SN��N���0�1�%�:�2�.�}���T�Ư�V��
�����!�u�4�6�w�5�W����Ƹ�V��Y��ʡ�0��%�<��2���Y����\��=N��Xʱ�u�=�&�<�w�����K�ƿ�]��C��ʼ�u�:�u�1�2�}�����Ƹ�VF��G��U���0�_�u�0��9��������9F��QN�����u�u�0�0�6�8�W���8����g��s8����u�u�%�:�2�.�$��������N�����;�u�u�u�>�}��������VN��Z��6���-�u�=�;�w�}�W�������e��S/�����,�i�u��#���������_��v
�����0�0�4�x�w�2����I���F�N��U���u�u�u�u�w�}�W���Y�ί�R��V��1���9�}��'�?�.�3��� ���r(��T*�����<��:��~�W�W���Y����Z ��N�����%�:�0�&�]�}�W�������Z��v
�� ���h�6�4�4�6�4�6�������X'��R�����9�,�d�n�w�8�Ϲ�����VF��Y/�����0��,�_�w���������V"��TךU���>�%�h�u�2�8����Y����w��a�����1��7�i�w���������C"�������&��9�,�f�}�9���=����R
��q��<��u�0�1�2�9�/��������V��R����_�u�x�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Y���a	��S��U���u�9�6�u�%�.����Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x��'�!�#�8�Ͽ�������TA�1���m��1��5�>����������TA�����u�;�_�w�p����V�ƪ�AF��N�����u�'�u�&�3�)�W���Y����F��V�����6�:�&�!�%�.�������K��V��ʳ�9�0�{�u�?�.�W���ӕ��E��XN�����9�u�0�4�w�5�W�������Z��_ךU����>�-�1�:�4�W�������G����U���&�8�9�1�>�}�����״�W	��^ �U���_�u�x��4�3�W����ƭ�VF��ON������a�u�:�9�8�����ƪ�AF����U���u�|�u��2�8�W��Y����F�������1�!�0�a�z�4�W���ӂ��]F��]����y�4�1�%�$�}��������F���U���d�u�:�4�9�W�W��Y���zF��CN�U���;�}�6�4�6�2���������C��4��� ��u�_�w�p�&ϱ����a	��SF��1�����1� ��}�W�������W��U'��\���x�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���T����X9��r�� ���!�4�%�<�0�4����Y����[	��h��1����u��!������0���K��X��ʶ�4�4� �u��)�1���+����9F������u��!��;�9�Ͻ�����_��X/��&���u��%� �'�)��������]��OT�����,�"�'�{�&�����*����Z��^ ������|�u�u�0�3�������9F�N��&���h�u��6�w�p�W���Y����T��E����!�u�c�o�w�W�W�������R�=N��U���4�%�0�9�w�}�W���*����V%��N��U���u�u�x�u�9�}��������F�N������>�-�u�j�}��������KJ�N��U���x�<�u�&�3�1����Y�����D�����u�u�k�6�2�8�2���Y���F�N�U���u�!�
�:�>�W�W���Y����R/��N��U��u��!���9����U���K�^ ��&���4�4�!�}��>�X��T�ƨ�D��^��U���u�6�4�4�6�4�>���D�Ư�R��V��!���1� �y�u�z�4�Wϭ�����ZǻN��U���!��!�u�w�}�IϽ�����\��B ��U���u�x�u� �w�(����������TC����!�u�|�u�w�}��������W)��S����4�4�<��#�f�W���Y����F��C
�����_�_�u�u�2�5��������	l�N�����&�6�4�4�%�0����P�����^ ךU���u��!��#�8���Yۉ��V��	F�����h�r�r�|�]�}�W����ƅ�Z������x�u�:�%�w�}�W�������|��R��<���h�6�4�4�%�0����Q����F�N��ʹ�:�n�u�u�2�9��������9F������!�u�i�u��)�8������]ǻN��1����!�u�i�w���������W�=N��U���!��!�u�k�}�3���6����^�UךU����!��!�w�a�W�������g��]����u��!��#�}�K���=����F��Z��\�ߊu�u��!��)�W��Y����R)��c��]���_�u�u��#�����E�Ư�R��B�����|�_�u�u��)�8���Y���P"��V!��!���}�|�_�u�w��������F��V�� ���8�}�|�_�w�}�3���6����Z�T*������8�}�|�]�}�W�������V�
N����� ��8�}�g�f�W�������|��N�U���!��!�0�'�l�^�ԜY�Ư�R��B�U��6�4�4� ��0�_��B�����C����i�u��!��)����H����F�T*�����d�u�h�6�6�<��������]ǻN��1����!�`�i�w���������W��d��U���;�u��n�