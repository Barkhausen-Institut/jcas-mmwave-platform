-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��GZ����x�u� �=�%�}��������K��E������:�0�!�w�������"��RT��Bʔ�2�&�u�e�b�p�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�U¶�u�e�`��'�/����7����]��~ �����;�&��'�8�<����T�ƍ�_F��P��U���0�#�1�x�w�<����ӯ��G��R ��U���0�;�9��1�/�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�x�u� �'�.�M��Y������G�����;�!�;�<�#�.�Ϛ�)���P	��^	�����:�u�u� �#�-�¿���� ��T������u�&�1�$�3����ӄ��P	��V�����<�=��y��q����*����@F��=C�U���u�;���2�W�������V��d�U���u�'�g��p�}�Ϝ�Q����W��@��Dʼ�u�<�&�u�9�>����Y����T��X�����<� �0�_�z�}�W���Y���F�N��U���u�u�u�u�w�>�������K�#���߇x�u���0�p�}��-����\��^�����6�;�7�u�2�4��������WF��E��ʡ�0��:�!�k�c�6���Y����]HǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�_�>�/��������F��RN�����!�
�:�<��l�C������F��^��[���0�<�
�!�y�1�L�������\��g�����4�9�9�4�;�W�Z��� ����@��C�����0�:�3�x��?����!����K%��R"��N��7�4�,� ���L��ӳ��`/��a�����;�&���]�p����������Y�����;�_�0�!�#�}����	����@F�N�����6�_�u�u��/�������F��^ �����4�u�h�3�;�8�}���Y����@��C��U���o�<�u�:�;�<�W������l�N������!��u�w�g��������]F�������n�u�%�'��}�Wϝ����	F����*���<�n�u�u�z�}��������GǻN��4���u�o�<�u�#�����&����\�N�����u�|�_�u�w�����Cӏ��@��[�����6�:�}�l�3�*����P���F��T��U��� �u�!�
�8�4�(������
F��@ ��U���_�u�u���}�MϷ�Y����_	��TUךU���x��!�_�w�}�5���Y����]F��S1�����#�6�:�}�`�9� ���Y����F�T,�����u�;�&�1�;�:��������Q��X����n�u�u�6�4�(�W����ƿ�W9��P�����:�}�b�1� �)�W���s���K��v-�� ���!�u�u�6�w�}�W����ƿ�W9��P�����:�}�b�1� �)�W���s���P6��YN��U���&�1�9�2�4�+����Q����\��XN�N���u�6�6� �w�}��������T��A�����b�1�"�!�w�t�}���Y����~6������9�2�6�|�]�3�W���=����lǑV�����!�'�u��w�;�2���
����ZǑN�����0�!�1�%�o�W�W�������PNǻN��U������u�w�}�W���Cӏ��V��T��D�ߊu�u�u����%���Y���F������u�h�d�_�w�}�W���>���F�N��U���u�;�0�0�w�`�F�ԜY���r3��e+��!���������W���Y�����[��U�����_�w�}�W���6����g9��c:��;�����
����Mϭ�����	[�z/��=��u�u�u����#���Y���F�N�����u�h�w���	�L���Y����p'��e+��U���u�u�u�o�>�)����C����9F�N��'���u�u�u�u�w�}�W������V�
N����u�u�
���}�W���Y���\��C����u����u�W�W���Y����j/��r)��U���u�u�u�;�2�8�W��H���F�t/��,������u�w�}�W�������	[�d��U�����u�u�w�}�W���Y����Z��P��O���n�u�u�u���W���Y���F�N����#�6�:�u�j��D���?����u ��d��U�����u�u�w�}�W���Y����Z��P��O���n�u�u�u���4��� ����tF�N����2�'�o�u�l�}�W���6����v4��N��U���u�o�<�!�0�/�M���B���F��v:��'���u�u�u�u�w�g��������AF��6��E��e�e�e�e�l�}�W���)����F�N��U���u�o�<�!�0�/�M���B���F��r"��4���u�u�u�u�w�g��������D��d%�����u�u��
��	�%���Y���\��C����u�����f�W���Yӵ��l4��y*��2����u�o�&�%�3�W��[����~'��UךU���u��
���}�W���Y�����^ ��O�����w�_�w�}�W���&����F�N��U���u�!�<�2�m�}�:���&����F�N��0���������W�������\� ��%����w�_�u�w�}�$���0���F�N��U���!�<�2�o�w��2��P���F��E��U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u��}�W���Y���F��^ �����9�2�6�#�4�2�_������\F��d��U�����u�u�w�}�W���Y���@��[�����6�:�}�l�3�*����P���F�v-��!���u�u�u�u�w�(�W���&����P9��T��]��1�"�!�u�~�W�W���Y���F�N��U���u�;�u�!��2��������W��S�����|�_�u�u�w��9���Y���F���U���
�:�<�
�2�)���Y����G	�UךU���u�� �u�w�}�W���CӉ����h�����0�!�'�d�w�2����I��ƹF�-��U���u�u�u�u�m�4�Wϭ�����Z��R����u�:�;�:�g�f�W���YӶ�F�N��U���o�:�!�&�3�1��������AN��
�����e�n�u�u�w��>���Y���F�N��Uʦ�1�9�2�6�!�>����Nӂ��]��G�U���u����w�}�W���Y�ƣ�GF��S1�����#�6�:�}�`�9� ���Y����F�N��'����u�u�u�w�}��������\��d��U������ �w�}�W���Y����@��[�����6�:�}�u�8�3���B���F��v<��6����u�u�o�>�}��������P]ǻN��U��������}�Mϱ�ӕ��l��P�����u�u����}�W���Y����]F��C
�����
�0�!�'�a�9� ���Y����F�N�� ����u�u�u�w�}��������T��A�����u�:�;�:�g�f�W���Yӥ��a?��d+��U���o�<�u�&�3�1��������AN��S�����|�_�u�u�w��#���7���F������ �:�<�n�w�}�Wϓ�5����})��N��Oʺ�!�&�1� �8�4�L���Y����e#��{!��U���u�o�:�!�$�9������ƹF�;��0����u�u�u�m�2�ϭ�����T��=N��U���������#������G��[���ߊu�u�u����3���:���	����*���2�6�_�u�w�}�2��Y���F�T�����!�
�9�2�4�W�W���Y����F�N��U���u�;�u�!��1����s���F��v"��:���u�u�u�u�9�}��������l�N��6���u�u�u�u�w�}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u���W���Y���F��^ ����� �:�<�n�w�}�Wϝ�:����z(�N��Oʼ�u�&�1� �8�4�L���Y����v%��{N��U���u�o�<�u�$�9������ƹF�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U���� �����W������G��[���ߊu�u�u��w�}�W���Y�������*���2�6�_�u�w�}�$���Y���F�T�����!�
�9�2�4�W�W���Y����*��e<��;���u�;�u�!��1����s���F��c/��8���u�u�u�u�9�}��������l�N��'���u�u�u�u�w�}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u��	�#���Y���F��^ ����� �:�<�n�w�}�Wό�-���F�N��Oʼ�u�&�1� �8�4�L���Y����`2��N��U���u�o�<�u�$�9��������F��SN�����0�!�_�u�4�3����Y����U5��E��Oʦ�'�;�u�h��)���*����VN��^��6���|�_�u�:�$�<�ϵ�����F��T�����2�o�u�0��-�O�������u��C*����u�6�;�!�9�}�9�������F��^ �����o�u�0��'�e����Q����@��C�����:�u��!�6�<����B���P	��C��U����1�u�u�w�}��������E��X��U���;�:�e�u�m�}�W���Y���F�N��U���u�u��!�$�i�8����Χ�Z��s��\�ߠu�&�2�4�w�}�2���Y���F��D�����6�o�u�e�l�W����s����v��R��R��"�0�u��:�/���Y������u#�����1�%�m�
�w�}�������V��^�����u�u�4�4�4�8�W���H���F��B�����u�k�e�_�w�}����D����F�N��U���u�u�u�u�w�}�W���Y���F�_��3ʺ�u�:�3�u�w�<����
����R��E �����!�h�u�4�$�q�W�������V��h�����
�0�0�!�8�)����G�ā�g%��d��Uʴ�<�%�!�h�w���������9F������2�h�u��:�/���Y����A��
P��;���'�2�y�u�w�}�W���Y���F�N��U���x�d�:�u�w��W���=����F�U1�����h�u��!��(���s���P��N�����k�e�_�u�w�<����
����TF�^�U���6�0�u�k�g�W�W������F��(��3�����w�_�w�}����D����9F������'�<�'�2�j�}�[���YӉ��\��R	��K��_�u�u�4�#�/�W�������V��^�E���u�u�%�0�w�c�F�ԜY�ƿ�_9��B �����4�>�h�u���:���[���F��[1�����k�w���{�}�Wϭ�����G��S�W�����w�_�w�}�������F��b"��&���u�u� �0�'�)��������GF�L��*�����y�u�w�(�������D��rZ�\��'�u�4�}�w�}����D�Ư�XJǻN��U��6�y�u�u�5�`�W���s���PF�F�����u�k�r�r�{�}�WϽ�����[�^�����u�6�;�h�w����Y����P��
P��7���y�u�u�%�>�}�IϽ�����F�T�����6�;�h�u�g�q�W�������Z��YN��U��y�u�u�4�8�)�J���8����l�N�����h�u��:�#�W�W�������R��B��Kʺ�0�y�u�u�:�1�������F��R �U���%�h�u��]�}�W�������W��T��Kʺ�0�y�u�u�'�)��������[�X��Y���u�:�0�3�8�}�Iϱ���ƹF��Y
�����u�k�:�0�{�}�WϽ�����GF����ߊu�u�6� �w�c������ƹF��G����u���1�{�}�WϿ�����[�^�E���u�u�6�'�.�3����G����D�N�����u�k�r�r�]�}�W���K���P#��N�U��<�u�&�1�>�}����HӠ��\��=N��U���9�8�1�u�i�z�P�ԜY�Ư�QW�	N����_�u�u�0�e�`�W���;����F�T��H���d�y�u�u�4�>�������W�=N��U���u�k�6�;��q�W�������_F�I�Y���u�6�%�h�w��5���s���P��[�����;�h�u�d�{�}�WϬ����A��d��Uʧ�!�9�8�1�w�c�P���s���A��S�R��_�u�u�&�4�`�W��U�����V�����<�u�k�r�p�W�W���
���F�BךU���&�6�'�u�i�z�P�ԜY�ƾ�G�	N��R��u�u�_�;�w�	�L�