-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B6��V�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mώ�0����KǶN����g�u� � �#�o�F�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�}�|�g�f�}��������}��X ��U���!� �0�!�w�2��������K��[�����&��&�'�2�W�Zϐ�����_F��D�����&��!�'�6�}��������]l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z��������2����������6�:�2����Yӯ��F��V ��:��� �&�4�0�<�-�W�������@��V��U���x�u�=�u�6�-����Y����Z�'�����9�,�!�0�2�<�ϸ��Ɗ�aF��[��ʼ�%�0�0�!�3�p�W���Ӎ��^%��Q>��%���0�>�%�z�w�2����������(��[���_�x�u�u�w�}�W��T���K�C�X���u�u�x�x�]�p�>Ϸ�Y���OF��eN�]���;�<�0�u�z�p�W���T���K�������u�u�u�)�w�p�Z��T���K�C�U���x�x�_�x�w�}�WϢ�Y���K�C�X���x�x�u�u�+�p�W���Y�����~<��U�6�:�&�u�+�p�W���T���F�N��U���x�x�x�x�z�p�Z��T���OF�Kd�U���u�u�u�u�w�}�W���Y���F�N��U���u�_�x�u�w�}�W���T���K�C�X���x�u�u�)�w�!�Z���Y���K��(��U����6�:�&�w�!�Z��Y�ư�K�N��U���x�x�x�x�z�p�Z��T���F�N�����u�u�u�)�w�p�Z��T���K�C�U���u�u�x�x�]�p�&Ϸ�Y���OF��eN�]���;�<�0�u�z�p�Z���Y�ư�K�������u�u�u�u�w�p�Z��T���K�C�U���u�u�x�x�]�p�Z�������]��R��O���u�u�=�u�>�8����������VN�����:�u�3�>�'�}����7����V ��E>���߇x�u�u��3�/����s���F�N��6���_�x�u�u�w�}�'��K���F�V��%��a�x�u�u�w�k�$���Y���9K�N�����;�u�0�4�m�p�W����ƭ���YN�����u�3�6�0�1�>����C����(��t��%���=�&�~�1�2����s��� �������;�8�0�u�1�>��������@\�_�;���:�3�0��6�8�6�������TǶd�U���3�<�<�;�w�2�ϑ�����K�-�����<�;�&�4�2�1����Y����G����ʡ�0�=�2�0�#�4����Y����Y��^ ��X���u�:�;�7�w�����
����R��C��Yʸ�1�}�z��:�2���Y����G��`�����u�u�-�8�;�}����Y����RF��R�����&�u�4�0�]�p�Z���Y����
��S��U���u�:�3�<�>�3��������@��C�����3�0�u�:�#�8��������GǶN�����0�{�u�=�9�.�Ͻ�����]F��C��6����h�d�{�w�5����
ӈ��]����U���6�&�x�u�w�8� ���Y����P	��Q�����{�u��0� �}�����Ư�V��SN�����:�1�{�u��8� �ԑT����@F��R
��ʰ�4�9�u�u�?�;�W���������T�����&�!�0�6�2�;�����ƥ�G	��_חX�����m�&�w��W���Y������R��U���=�3�'�!�8�1�������\��^�����"�9�_�x�w�6��������]��Y
�����%�<�u�=�w�/����	����F�������:�1�y�!�2�9��ԑT����]F��X����� �<�2�!�2�1����7����V ��N��ʢ�0�u��0� �`�F���
ӓ��WF��Ed�U���=�u�:�3�>�4����s��ƴF�T-�����_�x�u�u�g�m�W�����ƴF�I�D���u�u�;�<�2�u�>�ԑT���V��N��<ʶ�:�&�u��~�p�W���^����[�������}��_�x�w�}�F��Y�Ɲ�Z��Y��$���x�_�x�8� �+�W�������@��V�����u��6�h�f�}�_�������V�d�Uʾ� ��0��%�5����Y���U��T�����0�!�u�:�6�t�Z���:����Z��Y������1�'�u�f�}�D���L���FǶN��U���u�u�u�u�w�}�W���Y����F��N�Y���y�x�u�u�w�}�W���Y���F�N��U��u�d�u�f�w�h�}��Y���F�N��U���u�u�u�u�e�q�E��H���JǶN��U���u�u�u�u�w�}�W���Y����F��N�Y���y�_�x�u�w�}�W���Y���F�N��U��y�d�y�d�{�}�[��Y���F�N��U���u�u�u�u�w�h�W��Y���W�=C�U���u�u�u�u�w�}�W���Y���R�X�U���u�_�x�u�>�8����=����[�N������>�6�6�2�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�Cװ���4�,�<�0�l�}��������@��[����c�{�9�n�w�(�Ϸ��Ȣ�^��T1��Ĵ�9�_�u�&�w�2��������A��R����_�;�<�,������������N�����6�_�u�u��>�W���Y���F������u�4�2�u�w�2�F���D����9F������3�0��4�2�g��������R��\����u�h�a�|�]�}����s���`��[�����u�u�u�u�9�.��������F�d�����>�-�u�u�w�}�ϭ�����Z��N�����0�u�u�u�w�}�W���ӕ��l
��^�U���6�:�3�0�w�}�W���Y�ƥ���h�����0�!�'�g�3�*����P���F��X�����u�u�u�u�w�3��������l��C��D���:�;�:�e�l�}�WϽ�����F�N��U��<�u�!�
�8�4�L�ԜY�Ư�R��Y'�U���u�u�u�;�$�9��������G	��Y�����:�e�n�u�w�>�������F�N����!�
�:�<��8����H�ƨ�D��^����u��!���}�W���Y����]F��S1�����#�6�:�}�`�9� ���Y����F�T*�����f�u�u�u�w�}�ϭ�����Z��R����u�:�;�:�g�f�W�������z��N��U���o�<�u�!��2��������W��S�����|�_�u�u��)�>���Y���F������9�2�6�#�4�2�_������\F��d��Uʶ�4�4�;�c�w�}�W���Y����G��X	��*���!�'�d�u�8�3���B�����C��<���u�u�u�o�>�}��������E��X��Bʱ�"�!�u�|�]�}�W�������F�N��U���;�&�1�9�0�>����������Y��E��u�u�6�4�6�3�N���Y���	F����*���<�
�0�!�%�l�W������]ǻN��1�����e�u�w�}�MϷ�Y����_	��T1�����}�b�1�"�#�}�^�ԜY�Ư�R��Y'�U���u�u�u�;�$�9��������G	��Y�����:�e�n�u�w�>��������F�N����!�
�:�<��8����H�ƨ�D��^����u��!���n�W���Y����]F��S1�����#�6�:�}�`�9� ���Y����F�T*�����d�u�u�u�w�}�ϭ�����Z��R����u�:�;�:�g�f�W�������z��N��U���o�<�u�!��2��������W��S�����|�_�u�u�4�<����I���F�N��U���
�:�<�
�2�)���Y����G	�UךU����!���w�}�W���Cӏ��@��[�����6�:�}�b�3�*����P���F��V����u�u�u�u�w�3��������l��C��D���:�;�:�e�l�}�WϽ�����bU�N��U��<�u�!�
�8�4�(������F��@ ��U���_�u�u��#��&���Y���\��YN�����2�6�#�6�8�u�@Ϻ�����O��N�����4�;�`�u�w�}�W���ӕ��l
��^�����'�d�u�:�9�2�G��Y����w��~ ��U���u�u�o�<�w�)�(�������P��_����!�u�|�_�w�}�3���0����F�N��U���&�1�9�2�4�+����Q����\��XN�N���u�6�4�4�9�e�W���Y����Z��C
�����
�0�!�'�f�}�������9F�������u�u�u�w�g��������T��A�����b�1�"�!�w�t�}���Y����R/��^��U���u�u�;�&�3�1��������AN��
�����e�n�u�u�4�<����H���F�N��U���
�:�<�
�2�)���Y����G	�UךU����!���e�}�W���Cӏ��@��[�����6�:�}�b�3�*����P���F��V����u�u�u�u�w�3��������l��C��D���:�;�:�e�l�}�WϽ�����bW��N��U��<�u�!�
�8�4�(������F��@ ��U���_�u�u��#��&��Y���\��YN�����2�6�#�6�8�u�@Ϻ�����O��=N��U���!��9�1�9�}�W���ƿ�W9��P�����u�6�4�4�"��W���Y����\��D�����6�#�6�:��m��������l�N����� ��u�u�w�}�W���Y����_	��T1�����}�e�1�"�#�}�^�ԜY�Ư�R��B��U���u�u�u� �w�)�(�������P��]����!�u�|�_�w�}�3���6����F�N��U���u�!�
�:�>���������W	��C��\�ߊu�u��!��)�C���Y���	����*���<�
�0�!�%�n�W������]ǻN��1����!�`�u�w�}�Mϱ�ӕ��l
��^�����'�f�u�:�9�2�G��Y����w��x��C���u�u�o�:�#�.��������V��EF�U���;�:�e�n�w�}��������F�N��Oʺ�!�&�1�9�0�>����������Y��E��u�u�6�4�6�(�>���Y���	F��CN�����2�6�#�6�8�u�GϺ�����O��N�����4� ��u�w�}�W����ƿ�W9��P�����:�}�e�1� �)�W���s���P"��V!��<��u�u�u�u�"�}��������E��X��Eʱ�"�!�u�|�]�}�W�������zW��N��U��� �u�!�
�8�4�(������F��@ ��U���_�u�u��#����Y���\��B�����:�<�
�0�#�/�D�������V�=N��U���!��!�d�w�}�W������G��X	��*���!�'�f�u�8�3���B�����C����u�u�u�o�8�)��������l��C��F���:�;�:�e�l�}�WϽ�����G/��N��U��:�!�&�1�;�:�������� V��X����n�_�u�u��)�8���I���F���U���
�:�<�
�2�)���Y����G	�UךU����!��!�f�}�W���CӉ����h�����0�!�'�f�w�2����I��ƹF��s��:���g�u�u�u�m�2�ϭ�����Z��R����u�:�;�:�g�f�W�������|��N��U���o�:�!�&�3�1��������AN��
�����e�n�u�u�4�<����(���F�N��ʦ�1�9�2�6�!�>����Iӂ��]��G�U���6�4�4� ��}�W���Y�ƣ�GF��S1�����#�6�:�}�g�9� ���Y����F�T*������u�u�u�w�}��������T��A�����e�1�"�!�w�t�}���Y����R)��fY��U���u�u� �u�#�����&����\�N�����u�|�_�u�w��������F�T�� ���!�
�:�<��8����J�ƨ�D��^����u��!��#�d�W���Y����F��C
�����
�0�!�'�d�}�������9F������!�d�u�u�w�g����
����\��h�����f�u�:�;�8�m�L���YӅ��G��C?�U���u�o�:�!�$�9��������G	��^�����:�e�n�u�w�>��������F�N����&�1�9�2�4�+����Q����\��XN�N���u�6�4�4�"��D���Y����\��D�����6�#�6�:��m��������l�N����� ��a�u�w�}�W���Y����_	��T1�����}�e�1�"�#�}�^�ԜY�Ư�R��B��@���u�u�u� �w�)�(�������P��]����!�u�|�_�w�}��������W)��N��Oʺ�!�&�1�9�0�>�}���YӅ��R��X�����u�o�:�!�$�9��������9��+�����9�9�:�n�]�<��������VF��{N��U���4�4�9�9�8�}��ԜY�˺�\	��D�����_�u�x�=�8��������P	��C��U���8�=�&�&�w�g�������F��G�N�ߊu�<�;�9�4�8�������\��C
�����u�h�r�r�]�}����Ӆ��@��[��U���u�!�
�:�>�}�J���^���@��V��'���!�:�;�u�w�}���������Y��E���h�}�!�0�$�c�G���s����Z��[N�����0�3�u�u�m�?�������U��RUךU���;�9�6�:�0�8����Y����\	��V ��Hʳ�9�0�_�u�>�3�Ͻ�����u ��[\��U���9�4�u�h�1�1��ԜY����R
��r �����0�u�u�u�8�1����DӀ��@��=N��Xʖ�0�_�u�<�9�1��������F�T�����:�<�
�}��0����
����\��XN�U��}�!�0�&�i�2����D����O��N�����u��0���}�W���Y����g	��E1������4�0�x�w�2����I����N��_��H���!�0�&�k�g�t�L���
����_F��X�����u�u�o��2�	�1���ۍ��^6��D��Dʱ�"�!�u�|�m�}�������\��E��R��|�_�u�<�9�1��������F�T�����:�<�
�}��0����
����\��XN�U��}�!�0�&�i�2����D����O��N�����u��0���$�W���Y����_	��T1�����}�u�:�;�8�m�W��Q����A�^��N�ߊu�x��!�]�}����Ӆ��G��~N��U���u�;� ��#��_������\F��T��]���0�&�k�:�?�/�J���^����F��P ��U���!���u�w�}�W�������R9��[�����:�e�u�h��)����Gۉ��V��	I�\��_�u�<�;�;�>��������C��N�����4�4�!�>�"�����T�ƨ�D��^��O���:�=�'�h��)����G���]ǻ�����6�4�4�:�%�(����Y����G"��V1������4�0�x�w�2����I����N��_��H���!�0�&�k�g�t�L�ԜY����R
��s��!���1� ��u�w�-�3���&�Χ�F��V��X���:�;�:�e�w�`�_������	��R��K��|�n�u�&�0�<�W�������W��U'��Oʆ�6�4�4�!�<�(�'�������W	��C��\��u�:�=�'�j�u����
���O�=N�����9�6�4�4�8�9�$���:����C��C��]���8�=�&�&�f�9� ���Y���F��C����:�=�'�h�p�z�^�ԜY����R
��s��!���1� ��u�w�-�3���&�Χ�F��V��X���:�;�:�e�w�`�_������	��R��K��|�n�_�u�>�3�Ͻ�����\��B ��U��� �%�!�4�6�)����T�ƨ�D��^��O���:�=�'�h��)����G���]ǻ�����6�4�4�'�:�2����Cө��C��V��¾�%�x�u�:�9�2�G���D�Σ�[��
P�����&�k�e�|�l�W�W�������w��x�����u�u�u� �'�)��������W	��C��\��u�:�=�'�j�u����
���O�=N�����9�6�4�4�"�	����Y����F��C*�����d�u�:�;�8�m�W��Q����A������k�e�|�n�]�}�Zϊ�����V
��DN��ʼ�u�4�%�0�;�o�W������P	��C��U���%�!�0�4�w�}�W�������AF��]�X���-�'�u��1�/����ZӅ��UF��T�����3�'�<�u��/����=����9F��X �����>�<��4�2�8����Cӏ��V��T��2���=�&��0����������[��N��F�ߊu�:�&�4�#�6����-����V
��T�����0�u�h��#�9��������R��y�����&�>� ��2�����
����F��Y������1� ��;�$�W���Y����T��S��N���6�;�!�;�w���������JF�N�����'�o�u�n�]�}�ZϚ�����Q������!�0�1�9�.�4�W���	����XF��T��Uʶ�;�!�;�u��)�!�������\��Y�����h�}��%�#�8����Y����c��R*�����u��1�'�%�8����s���F�N��U���u�u�u�u�w�}�W���Y���F�������9�,�~�<�2����=����I��=d�����4�u��!��1����=���\��C
�����
�0�!�'�<�4�'�������JK��S�����|�o�u�:�?�/�J���^��ƹ��Y�����4�4�<��3�/����Y����_	��T1�����}��1�'�%�8����Y����G	�N�Uº�=�'�h�r�p�f�}���������C�����'�8�;�u�m�.�������F�UךU���;�9�6�4�6�<����8����QF��D�����6�o�u�e�l�}�����Ư�R��V��!���:�%�u�u�#�����Y���A��=N�����7�!�u�0�'�g������ƹ��E�����0�%�:�u��<�������F�N����4�u�&�w�%�8�L�������Q����*���:�!�u�;�2�8�L�������Q����*���:�!�:�u��<�������	F��P ��U���d�n�_�0�>�W�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d��X���'�4�0�4�w�3����
����_F��EN�����2�!�0�1�#�}�������KF����Uح�6�:�>�u�z�}�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�'�4�2�3�������C��R��&���9��>�_�w�8��ԜY�ƥ���^ �����}�4�%�0�;�t����s���F��X	�����i�u�:�u��:����B����������;�u�'�6�$�f�}�������v��[��O���%�:�0�&��0�������F��P��U���<�u�<�<�0�8��������p
��OG�����u�u�u�6�8�:�������F��X	�����_�u�u�u��:����=����[��c������9�_�u�w�}�2�������AF�S��!���9���9�w�2�W�������U"��d��Uʰ�1�<�n�u�2�9��������9l�C��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�2��������	��^ ��6��� �!�u�x�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F��\�����:�3�<�<�9�.����������U�����=�u�9�d�w�2����Y����G��D�����x�u�=�8�#�}�����Դ�W	��^ �U���u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W�������VF��G-�����%�<�2�u��-��������]�������"�'�{�$��8�$�������4��d��Uʲ�;�'�6�8�'�u�W���YӍ��^6��D��U���u�h�u��:�5����Y���F�N��Uʼ�!�2�'�'�9�8�FϪ�Y����RǻN��U���8�:�3�0��<���Y����p	��g�����|�u�x�<�w�4����Ӕ��T���A���h�m�u�u�'�/�W���Y���F�d�����>�u�h�u�6�-����U���K��YN�����:�<�_�u�w�}��������KF�=�����9�g�y�u�z�4�Wϭ�����ZǻN��U���4�9��0�w�c��������V�C����7�:�0�;�w�}�WϽ�����_F�S����3�0�y�u�w�p�W���Y����_	��T1�����}�u�:�;�8�m�}���Y�Ư�\��^ ��U��u��0��9�}�W���Tӏ����h�����0�!�'�d�w�2����I���F�T-�����u�u�h�u��8� ��Y���K��YN�����:�<�_�u�w�}�4���-����F�������y�u�u�z�2�ϝ�����Z�������&�&�d�1� �)�W���Y�����R��<���u�k�6�:�1�2�4���Y���\��t��!���'�!�>� ��<���Y����G	�d��U���6�:�3�:��}�J���:����\7��N��X��� �u�:�3�8�4�(���7����R��_�����:�e�_�u�w�}�4���-����F�������y�u�u�z�2�ϝ�����Z�������&�&�d�1� �)�W���Y�����R��4���u�k�6�:�1�8����Y���\��D�����6�#�6�:��}�������9lǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z���������@�������_�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԜY����[��N�����6�u�u�<�>�:����Y����V��N�����'�u�0�1�w�2�W����ƭ�Wl�C�����e�&�!�'�"�5��������AF��EN����4�4�<��'�}����
Ӓ��R��B �����u�x�u�=�w�4����ӂ��R���U��� �u�0�4�w�;����?���F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�0�2���������F��X���8�9��>�]�}����s���Z ��^�����2�}�4�%�2�1�^Ϫ����F�T<�����,�i�u��$�)�}���Y�ƥ���D��R��4�1�6�0�2�����^Ӓ��]l�N��Uʶ�0�0�� �#�a�W�������]��\��1����9�1�<�2�v�[���
����F��[�����_�u�u�u�w��������A��d��U���0�&�3�6�2�8�4�������[��N��U���6�0�0��"�)�K�������V��e�����;�x�|�_�w�}�W���+����v��S��D��u�u�u�0�$�W�W���Y�Ư�V��r��I���e�n�u�u�w�8�Ϸ�B����������;�u�'�6�$�f�}���+����u	��Y��U��;�!�6�0�2���ԶY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x��!�u�9�(�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d��X���0�=�%�u�?�}��������R��N�����4�&�;�u�8�)�ϛ�	����_��EךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z����Ƹ�VF��G�����u�:�4�u�%�<�Y�������`��D�����"�9�u�6�"�1�ϼ�Y����l�T*�����}�|�u�h�4�<����I���P"��V'��]���u�h�6�4�6�3�F�ԜY����R/��\��U��6�4�4�;�e�W�W�������U�R�����4�;�f�_�w�����0���Z�T*�����a�_�u��#��>��Y���P"��V'��@�ߊu��!���k�W��Y����R/��UךU���!���b�w�a�W�������]ǻ������m�u�i�w�����0��ƹ��C��<��u�i�u��#��>��YӅ��G��~F�\��u��!���m�}���=����]/�G��Hʶ�4�4�;�d�l�}��������T�S��1�����g�_�w�����0����Z�T*�����d�n�u�6�6�<����M�����C��<��_�u��!���F���E�Ư�R��Y'�N�ߊu��!���m�W��Y����R/��UךU���!���d�w�a�W�������]ǻ������g�u�i�w�����(��ƹ��C��$��u�i�u��#��&��YӅ��G��fF�U��u��!���f�WϽ�����bN��N�U���!���n�w�>��������F�������n�u�6�6�<����P�����C��$��u�6�4�4�9�u�^���DӅ��G��fV�Uʶ�4�4�;�}�~�}�JϽ�����b_��N�����;�}�e�u�j�>��������9F��s��<���d�|�i�u��)�>���H���P"��V'��]��u�h�6�4�6�3�F��YӅ��G��fF�\��u��!���n�}���=����]7�G��Hʶ�4�4�;�d�l�}��������S�S��1�����`�_�]�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǻC�<���!�&�8�9�9�}������ƹK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�x�u�z�W�W��Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x�#�:�>�2���������C
��PN�����4�%�0�-�w�p��������w��~ ��1�����>�%�z�}�������F�A�����6�4�4� �w�����>����@/ǻC�����
�u��!��1����Y����R0��^
�����_�u�;� ��0����CӃ��Z��@��[����%�!�4�'�4����-��ƹF��R �����4�u�_�u�w�}�$���Y���F�N��Kʾ�%�y�u�u�w�}�W���Y����]F��Y�����4�2�u�u�8�l�W��A���F��y�����0��4�0�j�}�9�������A6��D��U���<�u�<�!�0�/��������\F��T��M���u�%�'�u�6�}�}���Y�Ɵ�^��t��U���u�u�u�k��0�������F�N��U���u�u�x�<�w�.������ƹF�=�����9�g�u�u�w�}�J�������p
��OB��U���u�u�u�u�w�p�W���Y����_	��Td��U���6�0�0��#�}�W���Y�����D�����u�u�u�u�w�}�W���Y����]F��C
�����_�u�u�u��<�������F�S����7�0�3�'�w�}�W���Y���F�N��Uʷ�:�0�;�u�w�}�������F�N��U��u��!���6���Y����G	�B��X���;�u�;� ��)�(���*�����Y�����u�u��!��)�W���Y���[�T*�����'� �&�y�w�}�W���Y���F��CN�����4�4�!�}��>�X��T�ƨ�F�N�����4�<��u�w�}�W�������e��S'��U���u�u�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u��!��;�9�������F��V�������:�%�{�}�W���Y���\��D�����6�u�u�u�4�<��������F�N��U���!��9�1�%�0���Y���F�C�� ���!�
�:�<�]�W�W�������VF��G'�� ���8�9�;�u�9�(�$�������F�A�����6�4�4�;�4�<����Q����W��X����_�u�x�=�8��W���������C��2���%��u�x�!�2��������e��S:�����&�:�0�_�w�p����&�Ư�R��V��:���:�0�_�u�9�(�$���������^�����{�$��%�#�<�����Ξ�OǻN�����<�u�4�u�]�}�W���*���F�N��U���k�>�%�y�w�}�W���Y���K��YN�����0�u�4�2�w�}���Y���9F�N��;���:�3�0��6�8�J���7����V ��E>�����u�x�<�u�>�)��������T��XN�U��m�u�u�%�%�}����s���F��Z��6���u�u�u�u�w�c�$�������F�N��U���u�u�u�u�z�4�Wϭ�����ZǻN��U���%�0�9�g�w�}�W���D�Ɵ�^��t�����u�u�u�u�w�}�W��Y���@��[�����u�u�6�0�2�����Y���F������-�y�u�u�w�}�W���Y���K��YN�����:�<�_�u�w�}�2�������AF�N��U��6�;�7�0�1�/�W���Y���F�N��Xʼ�u�7�:�0�9�}�W�������z�N��U���u�h�u��#��&ǵ�	����W	��C��\���x�u�;�u�9�(�3���&�Χ�C�
�����_�u�u�u��)�8���Y���F�S����4�:�'� �$�q�W���Y���F�N��ʜ�%�!�4�4�#�u�$���V���F��N��Uʶ�4�4�4�<��}�W���Y����w��a�����u�u�u�u�w�}�W���Tӏ����h���ߊu�u�u��#���������C�	N�����u�u�u�u�w�}�W���Y���K�X�����9�2�6�u�w�}��������W)��N��U��u�%�;�n�w�}�W���Y���F�N��X��� �u�!�
�8�4�}�ԶY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x�� �u�:�)����?����Z
��EךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǻC�<ʜ�9�;�u��w�/����Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x��&�4�#�<�ϵ�	����v��^�����6�8�:�0�#�q����Y����R��Y	��;���=�&�&�u�z�}�Ϙ�+Ӗ��@��N��ʾ�%�z�u� �'�)�W���Y����J��E�����_�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԜY����Z��X��<��u�3�'��>�}�W�������[��DC����'�!�_�u�w�p����&�Ɖ�C ��p��ʐ�%�<��:�'��}���Y�˺�\	��VN������8��u�w�p��������_��V�����g�_�u�u�z�5����Y����U/��T-������u�u�x�!�2��������d��t��"���,�e�_�u�w�p����&�Ư�R��YN�����:�'� �&�]�}�W�������RF��V������u��!��1��������9F�C�����
�u��!�"�}�3���-����`��~F�����u�-��'�%�(�>���Y����G��X��0���<��:�%��	�^���Y����V��^�����_�u�u�u�w�����
���F�S�����4�0�y�w�}�W���Tӏ����R	��U���2�u�u�:�o�g�W�ԜY���F��B�����'�=�&�u�i�6��������c��RB��X���;�u�;�0�2�}����Y�Ƹ�R��S�����u�u�u��8�-����Y���[�~G��U���u�u�u�u�w�}�ZϷ�Yӏ��V�������u�:�b�o�w�W�W���Y������FךU���u�u�9�u�w�}�W���D�Ɵ�^��t�����u�u�u�u�z�4�Wϭ�����ZǻN��U����!��u�w�}�J���=����\!��B��Y���u�u�x�<�w�����������Z>�����d�1�"�!�w�t�W���Y����w��a�����h�u��!��1��������F�N��Uʦ�1�9�2�6�w�}�W�������z�N��H����0���{�}�W���Y���F��N������'�!�u�w�}�WϽ�����F�N��U���0���,�g�q�W���Y���Z�D�����6�u�u�u�w�>�������F�������1� ���t�L��Y����@��[�����6�:�}�b�3�*����P����]��R ������;�<��8�-�>��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�u�'�$�}�>�������9F�N�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x��.��������`��N������:�%�6�:�2����UӃ��[F��Y�����u��8�=�$�.�W��Y����z4��_������0�>�%�x�}�����ƭ�VF��CN��ʧ� �1�1�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F��Y(��2���%��o�u�1�/�>Ϸ�Y�Ƹ���Z>�����d�2�;�'�#�W�W���T����X9��r�����:�%��%�>�����:���F�A�����>�'� ��:��W���Tސ��\��-��U���%�0�9�g�]�}�W�������RF��X��ʶ�:�3�:��w�}�Z¨�������R��U���0���,�f�W�W���T����X9��T*�����6�4�4�:�%�(��ԜY���E��\1�����4�4�<��w���������t��GךU���x�=�:�
�w�����Y����R2��S
������_�u�u�&���������	F��C��U���>��%�<��2����-��ƹF�	�����u�4�u�_�w�}�W���7����R��N��U���k�>� ��6�8�[���Y���K��YN�����0�u�4�2�w�}���C����F�N������0��'�?�.�W�������\��R�����u�x�u�;�w�3����Y����VF��C��M��u�_�u�u�w�}�0���	����F�N��Kʜ�u�u�u�u�w�}�W���Y����]F��Y�����4�2�u�u�8�j�M���s���F��E�����_�u�u�u�w�1�W���Y���[�d�����>�-�u�u�w�}�W������G��X	�����u�u�u��#��W���Y���P"��V:�����&�y�u�u�w�p����0����w��h��;���=�&�&�d�3�*����P���F������9�1�;�h�w���������t��G�U���<�u�&�1�;�:����Y�����R��U���u�h�u��2�	�>��Y���F�C�����0���%�)�W���Y����p	��`��U���h�u��0� ����U���F�N��Uʦ�1�9�2�6�w�}�W�������F�N��H����!���3�(�>���P���F��CN�����2�6�#�6�8�u�@Ϻ�����Oǻ��U���0�4�0��9�4�0���	����9l�C��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�}����Y����t��GךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Zϗ�
����Z�������%�<��8�-��������@J��V�����4�;�;�u��0����
���F��(��U���&�&�u��2�6���Y����F��V�����,�!�'� �3�9�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d��2���<��:�%��g�Wϸ�ӯ��]F��C��;���=�&�&�d�0�3����s���K��X��ʐ�%�<��:�'�����>����b%��N��Xǣ�:�>�4�>�%�(�9���0���K��_��*���9�u�4�%�2�1�E�ԜY���E��\1�����3�;�6�:�1�2�4���Y����[	��h��6����u��0� ����s���K��X��ʶ�4�4�;�6�6�<��������F�C�����4�6�4�4�6�4�>���=����R
��c�����_�u�u�x�?�2�(���6����GF��V������7���]�}�W���?����\��t����!�u�:�>��-�������a2��=N��U���0�0�<�u�6�}�}���Y���X(��g�����u�u�u�k�<�(�'������F�N�U���u�;�0�0�w�<����Y���\�d��U���u�>� ��2�����
�����Z-������4�0�u�z�}��������AF��Y	��Gʡ�u�m�o�u�]�}�W���Y����F��ZN��U���u�k��u�w�}�W���Y���F���U���0�0�u�4�0�}�W���N���l�N�����u�4�u�_�w�}�W������F�N��Kʆ�8�9��>�/�}�W���Y�������*���<�_�u�u�w�}�3���0���F�	N�����:�'� �&�{�}�W���Tӏ��/��B�����}��8�=�$�.�FϺ�����OǻN��U����!��9�3�3�J���=����R
��c�����y�u�x�<�w�.������ƹF�N��6����u�u�u�j�}�4���-����F�N��U���x�<�u��2�	�1������F������u�u�u�h�w�����8���J�N��U���<�u�&�1�;�:����Y�����C��U���u�h�u��#�	�6�������zO�C����&�1�9�2�4�+����Q����\��XN����;�u�0�0�6�8�0�������F��tUװU���u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�}�Z���Y����]��~<�����&�u�x�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Y���z��V �����>�%�z�u�&������Ư�^��R ��Yʰ�6�u�:�!�>�4�ϵ�����@��N�U�����%�4�2�s�W���Y����T��B�����'�u�:�u�2�}������ƹK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�0��%�/����0���U	��~N��U���:�>� ��6�8�Z�������GǻN��X���:�
�u�$��/����Y����Z��X��<�ߊu�u�x�=�8��W�������^F��N��Xǣ�:�>�4��<�����:����9F�C�����
�u��0��}�4���-����F�C�����4�6�:�3�2�>�������� OǻN��X���:�
�u��#��W�������A	��D?ךU���x�=�:�
�w�����������C�����:�'� �&�w�}�Z¨�������C��U���!���1�"��_���Y����B��E)�� ���-�u�;�<�.�*��������t��GN��!���u�u�u�2�9�/�ϳ�	��ƹF�N��;���=�&�&�u�w�}�J���7����R��N��U���u�x�<�u�>�)��������W��XN�O���_�u�u�u�w���������[��S�����0��'�?�.�[���Tӏ����R	��U���2�u�u�:�c�}�J��Y���F��p�����u�u�u�u�j�}�^���Y���F�N��U���<�u�<�!�0�/��������\F��S�����u�u�:�!�:�-�_���Y���%��N��U���u�h�u�4�'�8����U���F�C����&�1�9�2�4�}�W���YӅ��G��N��U��u��!���2����Y���K�^ ��<���!�4�4�!�<�(�'�������W	��C��\���u�u�u�6�6�<����0�����C�����:�'� �&�w�p�W���Y����_	��Td��U���u�6�:�3�9�}�W���GӅ��V ��f'�U���u�u�u�x�w�3�W�������A9��N��U���6�:�3�0�w�}�W�������d��NF�Y���u�u�x�u�9�}��������F�N�����%�!�u�u�w�c��������W5��f'��\��x�u� �u�#�����&����\� N�����u�|�u�0�3�:�����Ƌ�] ��p�����n�_�u�x�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F��C�����u�:�8�!�?�����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�0�4�w�5�W���Ӑ��Z��^	��ʷ�u�=�u�4�2�-�����ƨ�_��V�����2�:�%�u�;�2�W��Y����G��S��U���<�u�'�8�#�8����Ӓ��G��X�� ���:�4�6� �#�;�Ϫ�Ӆ��PǻC����9�u�3�!�2��'Ͻ����v��^�����y�&�;�0�#�<�W�������]��R��[���x�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���=����R
��g��O���%�:�0�&��0�������F��P��U���<�u�<�<�0�8��������p
��OG�����u�u�u�<�w��������F��R ךU���u�u��!��1����=���F��C����e�|�_�u�w�}����Y����R0��^
�����h�d�u�=�9�}�W���YӅ��G��[�����,�i�u��#�����
������E>�����9�,�g�1� �)�W���_���F�N��U���u�u�u�u�w�}�W�������Z��X��N���u�u�0�1�>�f�W�������U]ǻ��U���6�&�n�_�w�p�����ƨ�_�������=�!�0�4�3�/����Y����W��_�����'�'� �&�w��ϱ����K��XN�����3�>�%�u�w�q����Ӓ��A��DN��ʴ�1�'�!�0�w�3��������F��D�Uʒ�;�1�0��2���ԜY����`��	N����'�!�_�u�w�9��������Z��=N��U���6�&�}�4�'�8����P�����^ ךU���u�3�'�&�9�����*����V%�������_�u�u�u�w���������W��[��Hʶ�4�4�4�<��9����Q����V��R�����d�1�"�!�w�t�Q���Y���F�N��U���u�u�u�u�w�}��������W"��s������4�0�0�6�p�^ϟ�=Ӆ��G��[�����;�n�u�u�w�8�Ϸ�B����������n�u�u�6�6�<����-����`��S��1����9�1�1�2��ǵ�����A��R��X���_�u�;�u�2�8����>����W��E����_�u�0��3�/��������F������2�;�'�!�]�}�W�������Z��v
�� ���h�6�4�4�6�4�3����Χ�Z��V�����x�|���4�<��������^/��=N�����0�0�4�0��3����-����_��=dךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Zό�����TF��SN�����6�:�&�;�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�����u�=�'�u�%�}�W���*���"��V����� �u�:�%�9�3����*��� ��'����u�x�u��4�o����(���g��RN��ʠ�0�u�:�4�3�2�W��������������0�8�u�;�#�8�W��Y����Z��^������0�0�4�$�}����Y����A	��E�����,�!�0�&�0�<�Ϸ�Y����F�-��G���:�4�;�&�w�5�Ϫ��Ư�]F�������u�;�!�0��6�Ϻ�����9F�d��X���0�:�1�!�2�8����KӞ��`��s=��Mʇ� �1�'�u�8�8����0�ƣ�VF��EN��[���=�&�_�u�z�<�ϫ��Ƹ���Y
�����m�7�!�1�#�}����������DB�����4�&�7�6�w�3����T�Ƹ�VF��\_�����<�{�u�x�]�}�Zϗ����F��B ��U���!���1�"��W���=����\'��d��6���u�x�u�u�"�}�Jό����P"��V:�����7��~�6�6�<����*����OǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z�+����ӣ��|��B�����;�_�u�x�?�2�(���=����]/��T*�����1��7��w�p��������w��~ ��U���!���1�"��}���T����X9��T*������6�4�4�8�9�$���:�����X��U���!���u��)�#�������zl�C�����4�6�4�4�"���������a	��S'ךU���=�:�
�u��)�8���Y����R ��Z<�����u�x�#�:�<�<��������W/��T*�����<���1�"�W�W���6����G5��G����0�!�!�u�8�6�2�������`��[��U��_�u�u�2�8�������F�N�����k�>�%�|�w�p��������V��V ��U���:�d�u�h�o�}�WϮ��ơ�CF�N��Uʆ�8�9��>�w�}�J�������p
��N��U���u�u�x�<�w�.������ƹF�=�����9�g�u�u�i�����:����F�N��U���u�;�u�!��2��ԜY���P4��R�����u�h�u��$�)���Y���F�C����&�1�9�2�4�}�W�������z��N��U��6�4�4�:�3�����Y���K��YN�����!�
�}�>�'�}�W���Hӂ��]��GךU���u��!���}�W���GӅ��G��v
�� ���y�u�u�x�w�3�W���=����GN��d��Z��x�u�:�;�8�m�}���Y�Ư�R��Y?��U���h�u��!������(���F�N��Uʆ�6�4�4�!�����K����W	��C��\���u�u�6�4�6�3�>���Y���P"��V:�����7��u�u�w�p����*����G��F�����u�|�d�1� �)�W���Y�����C�����;�u�k�6�6�<����-����`��N�U���u�!�
�:�>�W�W���Y����R)��~N��U��u��!��8�����U���K�X��:��� ��!�
���������\F��=N��U����!��!�w�}�W�������u��e�����u�u�x�u�"�}��������l��d��Dʱ�"�!�u�|�w�}�WϽ�����_��B��Kʶ�4�4�4�<��)�L���Y���	����*���<�_�u�u��.��������@\ǻN�����&�}��!��2�%�������w��q��'���1�|�u�u�5�:����Y����w��x�����u�h�}�!�2�.�IǱ�����A��G�U���u�6�4�4�"�	����E����G��DS����'�h�r�r�~�W�W���Y����zF��^��ʾ�%�x�u�:�'�}�W���YӅ��G��C:�����|�i�u��#���������zO��N��U���6�4�4� ��0�&Ǘ�Y����w��q��'���1�}�|�_�w�}�W���Y����l�N��ʥ�:�0�&�_�w�}��������F�
N����� ��8��g�f�W�������|��N��Hʶ�4�4� ��:��F��Y����w��x��G���h�6�4�4�"�	����K��ƹF��s��:���f�u�h�6�6�<�������]ǻN��1����!�a�u�j�>��������C/�UךU����!��!�b�}�JϽ�����G2��G'��\�ߊu�u��!��)�A���DӅ��G��C:�����|�_�u�u��)�8���N�����C�����%�}�|�_�w�}�3���6����F������!�0�%�}�~�W�W���=����F��N�U���!��!�0�'�u�^�ԜY�Ư�R��B��E��u��!��#�8����I��ƹF��s��:���d�u�h�6�6�<�������O��N�����4� ��g�k�}�3���6����^��\����u��!��#�l�W������|��R��]��n�u�u�6�6�<����M���P"��V!��!����d�|�_�w�}�3���6����F������!�0�%�}�b�f�}���Y����R)��f^��I����!��!�2�-�_���s���P"��V!��$���i�u��!��)����Q����F�T*������u�i�u��)�8�������O��N�����4� ��u�k�}�3���6����^��G�U���6�4�4� ��}�K���=����F��Z��A��u�u�6�4�6�(�&���E�Ư�R��B�����`�n�u�u�4�<����(���F��V�� ���8��c�n�w�}��������F�
N����� ��8��`�f�W�������|��N��Hʶ�4�4� ��:��O��Y����w��x��L���h�6�4�4�"�	����@��ƹF��s��:���d�u�h�6�6�<�������O��N�����4� ��d�k�}�3���6����^��_����u��!��#�l�W������|��R��]��n�u�u�6�6�<����J���P"��V!��!����d�|�_�w�}�3���6����F������!�0�%�}�c�f�W�������|��[��Hʶ�4�4� ��:��F���s��ƓV��e:��