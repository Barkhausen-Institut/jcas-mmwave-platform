-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��E>�����=�_�x��#�2�MϚ�Ӥ��VǶN�����4�u�'�?�4�g�'���&�޴�9K�s��O��u� � �!�e�l�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����}�|�g�d�w�2�����Ƃ�G��V����� �0�!�u�8�-�������'��<������&�'�0�]�p�9�������z��E������!�'�4�w�3��������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��/����s����[��T�����!�<�&�4�#�<����Y����]F��*��A���u�=�!�<�w���������[��=C����{�u�=�&�1�1��������J��[��3����9�0�u�%�5��������[	����X���<� �0�a�b�2�W���Y����^��gN��ʃ�'�0�x�u���W���ӡ��W�B	�Fĥ�3�{�x�_�z������ƈ�_��
N�� ���0��'�=�$�}�W�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠ9�7�4�,�>�8�L�������V��D�����6�d�c�{�;�f�Wϫ�ӏ��VH��Z�����1�4�9�_�w�.�W���ݶ��v��E�����9�n�_�;�>�$�2�������@��Dd�����'�6�_�u�w���������[��T�����0�u�4�2�w�}���Y���l�N������!��u�w�}�W�������	[��V��U��u�%�'�}�w�}�4���Y���F�N��U���
�:�<�n�w�}�������F�N��U���
�:�<�
�2�)���Y����G	�UךU����!��9�3�3�MϷ�Y����_	��TUךU����0��u�w�}�MϷ�Y����_	��T1�����}��0��3�5�FϺ�����O��N�����3�0�u�u�w�}�ϭ�����Z��N�����%�!�u�u�w�}��������T��A�����b�1�"�!�w�t�^����Ɖ�C ��g���ߠ_�'�=�!�4�(�ό�5Ӊ��v��^�����<�_�u�x�!�2��������Gl�C�����&�2�;�_�w�)����Y����p��Y1��Uʼ�u�'�4�u�<�(�4���)����R��N�����u�|�:�u�#�����&����\�N�����u�|�_�u�>�3�Ͻ�����R��N��U���3�=�<�
�w�`�_������	��R��K��|�n�_�u�.�8�WϚ�����Z��N��ʴ�'�,�}��:�2����)����W��X����u�3�&�1�;�:��������Q��X����n�u�&�2�6�}�3���:����F�N�����4�;�!�o�w�2����D�Σ�[��
P��R���_�u�&�2�6�}�6�������]F�N�����4�!�>� ��8�'�������F��@ ��U���o�u�:�=�%�`�_������V�UךU���;�9�6�1�2�����Y����C��C��]���8�:�3�0��<�������\F��T��]���0�&�k�:�?�/�J���^����F��P ��U���'�!�1�0��)�W���&����P9��T��]��1�"�!�u�~�W�W���������v
�����u�u�!�
�8�4�(������F��@ ��U���_�u�<�;�;�>��������I���*���<�
�0�!�%�o�W������F��F�����h�r�r�n�w�W�W�������p	��~ ������%�u�u�#�����&����\�N�����u�|�o�u�8�5���^���9F��^	��ʶ�4�4�;�<�2�}�W���Cӕ��l
��^�����'�d�u�:�9�2�G���D�Σ�[��S�R��n�u�&�2�6�}�3���/����z��G��Oʦ�1�9�2�6�m�}�G��Yӕ��]��T-�����<�0�u�u�w�g��������\�^�����u�4�!�<�"�8����Y�ƿ�A��d�����<� �0�>�2�}�Ͻ�����a��M�����u�<�;�9�>�}����[���R��^��ʾ�0�u�3�6�6�<��������Z��[N��Uȡ� �w�_�u�#�/����Y����	��T*�����<���%�w�}����ӏ����RL�Uʴ�!�<� �0�<�8�W�������d��G��U���;�9�<�u�#�(�U�Զ����9l�T-�����0�<�0�i�w�)�(�������P�������&�2�0�}��8�>���J���9F�N�����&��>�_�w�8��ԜY�ƥ���^ �����}�9�|�!�2�W�W���Y����U/��R�����0�i�u��2��%�����ƹF�������%�u�h�4�<����s���F��V�������%�u�j�>��������]]ǻN��U���0���%�w�`��������F�R ����u�0�1�%�8�8��ԶY����[	��h�����%�m��'�#�.�Cצ�Y����[	��h��3���!�:�3�!�"�W�W�������RF��^��1���u�'�0�u�z�+����Ӆ��P%��Q'�����0�<�0�u�z�+����Ӆ��Z�X����r�r�_�u�z�5����Y����F��t��6���;�e�_�u�z�5����Y������R��%���_�u�x�=�8��W�������z��GךU���=�:�
�u��4�WǱ�����A��d��Xǣ�:�>�4�6�4�(�W�������Z�d��Xǣ�:�>�4�6�9��W�������Z��g�����x�=�:�
�w�����
����V��Cd��Xǣ�:�>�4�6�4�3�_������V�=N��X���:�
�u��8�)��������Z�d��3���!�&�a�-�w�3��������v��D�U��_�u�u�2�8�������F�N������0�u�u�i�)���Y���F�C�����:�9�4�u�j�;����Y�����E�����u�h�u�'�2�}�W���Y���F��N�����;�o�u�4�$�W�W���Y����A��C��U��>�-�'��#��^���Tӏ����[��U��3�9�0�u�w�-�������F�N�����u�k��>�w�}�W���Y���F�N��Uʦ�1�9�2�6�w�}�WϽ�Y���X��t��<���&�/��%�{�}�ZϷ�Yӕ��l
��^�����'�g�u�:�9�2�G�ԜY���P'��YN��K���!�0�&�k�g�t�W���Y���Z�D�����6�#�6�:��d��������9F�N��4���!�h�u��2�����I���F�C�� ���!�
�:�<��8����K�ƨ�D��^��U���u�6�;�u�w�c��������C�N��U���x�<�u�&�3�1����Y�����N��H����!���'�q�W���Y�������*���<�
�0�!�%�l�W������l�N�����;�u�k�}�#�8����I���F�C����&�1�9�2�4�+����Q����\��XN����u�u��:�#�`�W�������Z�B��U���x�u� �u�#�����&����\� N�����u�|�u�u�w�>�W���Y����u��C/�����!�u�u�u�z�2�ϭ�����Z��R����u�:�;�:�g�W�W���Y����]F�	N�����&�k�e�|�w�}�W��Y���@��[�����6�:�}�b�3�*����P���F��g����u��1�'�?�4�_���Y���K��B�����:�<�
�0�#�/�C�������V�N��Uʶ�;��u�k�4�<��������Z��N��Xʼ�u�&�1�9�0�>�W�ԜY����F
��G�����0��4�0�]�}�ϵ�����U6��g����2�;�'�!�]�}�W���=����R��=N��U���u�u�;�e�#�}�9�������A6��D��U���0�4�0�u�w�}�Z¨�����#��s��M���u�u�x�#�8�6�ϵ�����\��Q�����u�u�x�#�8�6�ϵ�����R��Q�����u�u�x�#�8�6�ϵ�����R��QN�����u�u�u�x�!�2��������G��DS�E���u�u�u�x�!�2����������R������_�u�u�w�p����&�Ư�P	�������4�;��d�]�}�W���T����X9��T+��U���0��_�u�w�}�Z�������P$�X����r�r�_�u�w�}�Z�������P$��YN�����=�<�}�|�w�}�W������l��u��ʶ�4�4�=�<��v�^���Y�����X��U�����6�4�6�<����s���F�A�����6�u��1�%�(�_���Y���K��_��*����<�u��3�/����Q��ƹF�C�����
�u��:�#�>����:����/�d��U����%�&�a�/�}���� ӑ��XH��G*��A�����_�u�w�}�W�������^��d��U���u�u�>�<�$�����Y����R
��N��Xʼ�u�7�:�0�9�g�W���
���F�N�����&��!�u�w�c�������F��N�����;�o�u�4�$�W�W���Y���X#��E�����u�k�3�9�2�}�Z����Ʈ�\
��YN�U���&�_�u�u�w�}�������9F�N��U���9�u�u�h�w�1�[���Y���F�N��Xʼ�u�&�1�9�0�>�W���Y�����N��H���:�=�'�h�p�z�[���Y���Z�D�����6�#�6�:��d��������9F�N��U����<�u�h�w���������J�N��Xʼ�u�&�1�9�0�>����������Y��E�ߊu�u�u�u�w�����D�Ư�\��_��]���|�u�u�x�8�)��������l��C��G���:�;�:�e�]�}�W���Y�Ư�]'�S����3�0�u�u�w�}�W���Tӏ����h���ߊu�u�u�u�w��W���D����G��DS�E���u�u�u�x�>�}��������l��C��D���:�;�:�e�]�}�W���Y�Ư�P��S����4�=�<�}�~�}�W���Tӏ����h�����0�!�'�d�w�2����I���F�N����� �u�k�6�6�<����Q����F�C�� ���!�
�:�<��8����H�ƨ�D��^��U���u�u�u�6�w�}�W�������A)��'��U���u�x�u� �w�)�(�������P��Z����!�u�|�u�w�}�W�������F������=�<�}�|�w�}�Z����ƿ�W9��P�����:�}�b�1� �)�W���Y���F������h�u��1�%�5����R���K�X�����9�2�6�#�4�2�_������\F��=N��U���u�u����`�W�������Z��U��U���x�<�u�&�3�1����Y����]��R ������;�&��6�3�}���Y���F��V������!�i�u��9����Q����p	��g�����x�|�_�u�9�}��������F
��G�����0��4�0�]�}����	���F��V������!�"�0�w���������[��	_�����6�<�&��3�/���s����4��d