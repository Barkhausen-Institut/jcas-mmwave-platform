-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B��G�����<�2�#�1�z�}�����ƈ�]F��\��X���'�2�;�9��2����Y����lS��Od�U���0�u�u�0�#�0����I��ƴl�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�u�4�}�G��:����Z�� �����9��&�'�:�3�ϝ�����G��=C�4����2�!�u�2�8����T�Ƃ�G��V����� �0�!�u�9�8����0����^��X חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�Z�������V\ǶN�����:�%�;�;�w�<����ӂ��RF����U���%�0�9�u�8�<�Ͽ�Ӗ��@��^��ʡ�0�x�u�4�'�8����Y����Z�/��ʡ�0�<�%�!�3�)�W�������T��D��U���!�}�|�<�w�5�}������GF��C�U���&�8�!�=�$�)�ϒ�Y������E�����<�;�:�u��9���Y����K��B��ʱ�!�u�&�4�%�3��������[��^�����=�u�0�0�#�9���Y������E�����_�x�3�'�#�8�1�������A�CחXʅ�%�9�;�u�2�<�M��s����\��^�����:�1��1�%�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�Cװ���4�,�<�0�l�}��������@��[����c�{�9�n�w�(�Ϸ��Ȣ�^��T1��Ĵ�9�_�u�&�w�2��������A��R����_�;�<�,��-����*����Z��^ךU���0�<�}�u�w�6����Y���F�N��Oʼ�!�2�'�'�9�8�EϪ�Y���F��=N��U���8�:�3�0��<����Cӏ��V�������u�:�a�u�j�e�^�ԜY����l�N������>�u�u�w�}�W���ӕ��l
��^�U����8�9��<�%�W���Y����Z��C
�����n�u�u�6�2�8�2���Y���F�N��U���
�:�<�n�w�}��������V�N��U��<�u�:�9�6�f�}���Y����R/��N��U���u�u�u�;��-��������`��N�����u�|�_�u�w��������F�N��U���u�;� ��#��_ǵ�	����W��X����n�_�u�u��)�!������F�T��ʦ�1�9�2�6�]�}�W�������Z��p�����u� �u�!��2���Y����w��a�����u�u�u�o�8�)��������O��=��U����%�!�4�'�4��Զs����Z��C��U���u�3��%�9�(�$�������ZǑN����>�&�2�!�%�W�W�������@��Y
װUʶ�;�!�;�u��0����
�����R	��U��>�%�z�n�w�>�����Ƨ�E��B�����u�:�9�4�w�`�>����Χ�F��R�����&�|�_�u�$�:����=����] ��ON��U���;� ��!��u�$���Hӂ��]��G��H���!�0�&�k�8�5���^���l�D������!���e�}�W��0����w��h��;���=�&�&�d�3�*����P���	��R��Kº�=�'�h�r�p�t�}���������C��G���,�u�o��'�)����ۍ��^6��D��Dʱ�"�!�u�|�m�}�������\��E��R��|�_�u�&�0�<�W�������Z����U���
�:�<�u�j�z�P�ԜY����R
��s��#���1�3�-�o�$�9�������V�=N�����9�6�4�4�6�4�0���Y�ƿ�W9��P��O���e�n�u�&�0�<�W�������Z����U���
�:�<�u�j�z�P�ԶYӕ��]��T*������9�u�u�w�}�W��0����w��h�����z�|�d�1� �)�W���C����G��DS����'�h�r�r�~�W�W�������w��a�����'� �&�6�w�}��������	[�I�Uʦ�2�4�u��#���������F�N����9�2�6�o�w�m�L�ԜY����Z��RN�����u�!�<�2�]�}��������X�������4�4�<��e�}�Mϭ�����Z�C��W�ߊu�!�'�7�#�}��������	F��C���ߊu�!�'�7�#�}��������	��T*�����<��g�u�w�4��������9l��P�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W��=����z��CN��ʖ�:�>��:�$�3�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d��X���=�&�&�6�>�3��������[��Y��U���4�u�;�u�2�.����������^ �����!�_�u�x�w�p�W���Y����F��X�����<�&�u��$�4�W���Y����KF��Z��U���u�'�;�3�%�8�W�������F��ךU���<�u�=�u�;�o�W������F�=N��Xʁ�0�1�!�u�8�8�W�������P"��V'��E���&�!�0�:�3�.�W�������[��D�����4�&�_�u�z�/��������G��S��U���=�!�4�u�g�}�Ϫ�ӈ��@��V��Uʁ�<�u�&�'�&�4��ԜY����\��_��<���<�!�'�_�w�p�W��Y����GF��C��U��� �%�!��#�W�W��T���K�N��U���x�x�x�x�z�}�Z���Y���F�N��U���y�a�u�_�w�p�W���U���F�N��D���y�b�u�x�w�}�E���I���F�\�G���_�u�x�u�w�q�F���Y���K��_�@���x�u�u�a�w�o�W��Y���F��=N��X���u�y�d�_�w�p�W���U����F�=N��Xʅ�%�9�;�u�2�<�W���W�Ɵ�^��t�����:�&�}�u�6�-����K��ƹK��N�U���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�w�p�#���Y����GF�������u�=�u�;�"�}����Y����W	����U���9�"�;�u�"�>����s���K�e�����u�u�u�e�$�;�Ϻ��ƥ�9F�N�U���4��9�1�w�}��������[��V���ߊu�<�&��m�}��������R��R-��\���7�2�;�u�w�4�W�������W��d�����>�u�=�;�w�}�WϷ�Y����V��CS��Rʡ�0�_�u�u�w�}�3���0����KF�F�����h�}�!�0�$�c�G���B���F������9�1�3�-�k�}�G��Y���F��s��#���1�%�-�i�w�l�L��Y����_��_�����'�=�&�&�3�/��������F�N�����6�4�4�4�>��W��^����[��N��U���6�4�4�4�>��F���DӅ��G��[���ߊu�u�u�u��)�!�������Z�T*�����<��n�u�w�}����s���F�T*�����3�-�i�u��)�>���*�����Y��E��u�u�u�u�4�<��������KF������9�1�;�_�w�}�W���=����R
��p��U��6�4�4�4�>��L���Y����]��QUךU���;�u�3�_�w�3�W�������9l�C�����!�0�1�!�w�/�Ϫ��״�G	��_��ʶ�:�>�1�8�>�s�W�������C	��Cd��X���;�0�u�u�$�.��������_��CN���ߊu�u�x��%�)���*����R��N��X���9�d�u�u��6����Y���F��R ��U��e�u�_�u�w�p�FϪ�����X�N�U���x�u�u�=�9�k�J���U��ƹF�N����u�u�k�f�w�W�W�������	l�G������8�9��<�%�}�������F�^�����2�0�2�}�6�-����K����[��N��Uʳ�'��<�u�w�2����)����@K��[�����u�u�u�3�4�3��������[��N��U���u�6�4�4�9�;�Ǘ�Y����w��~ ��D���|�_�u�u�w�}����Y���F�������g�}�|�k�}�3���0����KN��\ ��%���0�|�_�u�w�}�W���Y����F�N��ʹ�:�n�u�u�w�>��������UT��S��1����9�1�3�/�W�W���Y����R0��^
��G���h�6�4�4�6�4�0���B����������;�u�'�6�$�f�}���TӴ��A��RN��ʱ�!�u�:�&�4�}��������V��DN��ʻ�"�&�u�4�6�}�#���Y��ƹK�E�����u�:�u�=�w�4�����ƣ�V��^�����=�'��o�w�-����
۵��C
��[��\���7�2�;�u�w�4�W�������W��d�����>�-�u�=�9�}�W���������N��U���8�=�&�&�f�1��ԜY���F��V��ح�9�}�|�i�w�����?�Դ�X(��g�����|�_�u�u�w�3�W���	���F��SN��N���0�1�%�:�2�.�}���T�Ɗ�AF����ʻ�8�0�u�3�4�8��������C��G�����0�'�4�2�w�3�W���	��ƹK�C�����u�;�u�4�6�+����Yӡ��v��x�� ��u�<�u�:�w�����������R�����u�x�u�0�%�<��ԜY�Ư�R��B����u�h�6�4�6�3�ݦ�I��ƹF��s��:���6�}��8�?�.�������\F��R�����4�;�-�9�l�W�W���=����R
��x�����h�6�4�4�6�4�1���B�����C�����:�'� �&�4�}�JϽ�����_��G\�����;�u�0�0�6�8�0�������G��dךU����'�4�u�3�}����Ӊ��P	��Q�����u�0�u�=�$�q�����Ʃ�G��q(���ߊu�x�!�0�w�8�����ƭ�WF��C��U���u�4�4�4�3�9��������F��^�����u��u�x�w�.��������U	��G�����9�2�8�;�w�5�ϩ�Y������Y	�����u�;�:�u�z�}��������p
��S�����!�!�0�0�3�}�#���Ӊ��G��(�����=�u�4�4�w�p�W���Ӈ��V��VN�����<�u�=�u�&�����
���G	��X�����0�3�'�!�2�}�Z����Ƣ�^����3���{�u� �u�#�.����Y����F�������;�u�:�%�#�4�}���Tӎ��VJ��XN��R���0�0�<�&�2�9��������#��q�����{�u��;�3�����C����UF��A�� ���0�u�0�0�6�8�W���<����|��QTךU���'�6�&�}�6�-����K��ƹF��R	�����u�u�3�'�$�3�(���۵��C
��[��\ʡ�0�_�u�u�w�}�Ͻ�����_��G\��R��!�0�_�u�w�}�W���TӴ��A��PךU���u�u�u��#�����Q���F��V�����-�e�n�u�w�}�W�������|��T��;���=�&�&�d�3�*����P���P"��V'�����n�u�u�u�w�8�Ϸ�B���F��Y
���ߊu�u�;�u�%�>���Y����w��a������9�i�u��)�!�������l�N�����4�<���8�-�;���E�Ư�R��V��2���n�u�0�1�0�3����Y����W��C��N�ߊu��!��#�a�W���������=N��Xʶ�4�4�4�<��)�����ƨ�G��V��U���!�2�!�u�2�<�����ƹ�V��X����� �%�!�u�4�<��������Z�T*�����<��!�6�l�}�Z���=����R
��c�����u�&�&�8�;�/����=����R
��x��U���u�9�:�<�w�/�Ϻ�����F������:�!�4�u�?�}��������C��Y
�����u�=�u�r�w�5����s�Ư�R��V��!���:�%�u�h�4�<��������A	��D"��N���;�u��n�